module odo_pre_mix(in, out);
    input [639:0] in;
    output [639:0] out;
    wire [63:0] total;
    assign total = 0 ^ in[63:0] ^ in[127:64] ^ in[191:128] ^ in[255:192] ^ in[319:256] ^ in[383:320] ^ in[447:384] ^ in[511:448] ^ in[575:512] ^ in[639:576];
    assign out[63:0] = in[63:0] ^ total ^ (total >> 32);
    assign out[127:64] = in[127:64] ^ total ^ (total >> 32);
    assign out[191:128] = in[191:128] ^ total ^ (total >> 32);
    assign out[255:192] = in[255:192] ^ total ^ (total >> 32);
    assign out[319:256] = in[319:256] ^ total ^ (total >> 32);
    assign out[383:320] = in[383:320] ^ total ^ (total >> 32);
    assign out[447:384] = in[447:384] ^ total ^ (total >> 32);
    assign out[511:448] = in[511:448] ^ total ^ (total >> 32);
    assign out[575:512] = in[575:512] ^ total ^ (total >> 32);
    assign out[639:576] = in[639:576] ^ total ^ (total >> 32);
endmodule

module odo_sbox_small0(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h04;
        mem[1] = 6'h16;
        mem[2] = 6'h19;
        mem[3] = 6'h2a;
        mem[4] = 6'h06;
        mem[5] = 6'h32;
        mem[6] = 6'h24;
        mem[7] = 6'h08;
        mem[8] = 6'h3d;
        mem[9] = 6'h0f;
        mem[10] = 6'h1f;
        mem[11] = 6'h0e;
        mem[12] = 6'h27;
        mem[13] = 6'h0d;
        mem[14] = 6'h14;
        mem[15] = 6'h0b;
        mem[16] = 6'h09;
        mem[17] = 6'h11;
        mem[18] = 6'h13;
        mem[19] = 6'h35;
        mem[20] = 6'h18;
        mem[21] = 6'h33;
        mem[22] = 6'h3e;
        mem[23] = 6'h2e;
        mem[24] = 6'h2f;
        mem[25] = 6'h31;
        mem[26] = 6'h28;
        mem[27] = 6'h2b;
        mem[28] = 6'h2c;
        mem[29] = 6'h0c;
        mem[30] = 6'h00;
        mem[31] = 6'h21;
        mem[32] = 6'h02;
        mem[33] = 6'h3c;
        mem[34] = 6'h2d;
        mem[35] = 6'h30;
        mem[36] = 6'h12;
        mem[37] = 6'h38;
        mem[38] = 6'h1e;
        mem[39] = 6'h26;
        mem[40] = 6'h22;
        mem[41] = 6'h03;
        mem[42] = 6'h1b;
        mem[43] = 6'h1a;
        mem[44] = 6'h01;
        mem[45] = 6'h37;
        mem[46] = 6'h15;
        mem[47] = 6'h0a;
        mem[48] = 6'h20;
        mem[49] = 6'h05;
        mem[50] = 6'h3a;
        mem[51] = 6'h3f;
        mem[52] = 6'h1d;
        mem[53] = 6'h3b;
        mem[54] = 6'h17;
        mem[55] = 6'h29;
        mem[56] = 6'h34;
        mem[57] = 6'h10;
        mem[58] = 6'h1c;
        mem[59] = 6'h23;
        mem[60] = 6'h25;
        mem[61] = 6'h07;
        mem[62] = 6'h36;
        mem[63] = 6'h39;
    end
endmodule

module odo_sbox_small1(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3a;
        mem[1] = 6'h11;
        mem[2] = 6'h3d;
        mem[3] = 6'h00;
        mem[4] = 6'h32;
        mem[5] = 6'h37;
        mem[6] = 6'h15;
        mem[7] = 6'h1a;
        mem[8] = 6'h3e;
        mem[9] = 6'h33;
        mem[10] = 6'h3f;
        mem[11] = 6'h2b;
        mem[12] = 6'h19;
        mem[13] = 6'h0b;
        mem[14] = 6'h09;
        mem[15] = 6'h24;
        mem[16] = 6'h29;
        mem[17] = 6'h20;
        mem[18] = 6'h25;
        mem[19] = 6'h39;
        mem[20] = 6'h13;
        mem[21] = 6'h1d;
        mem[22] = 6'h26;
        mem[23] = 6'h34;
        mem[24] = 6'h10;
        mem[25] = 6'h2f;
        mem[26] = 6'h08;
        mem[27] = 6'h06;
        mem[28] = 6'h01;
        mem[29] = 6'h23;
        mem[30] = 6'h38;
        mem[31] = 6'h0a;
        mem[32] = 6'h2a;
        mem[33] = 6'h1e;
        mem[34] = 6'h03;
        mem[35] = 6'h22;
        mem[36] = 6'h2c;
        mem[37] = 6'h0d;
        mem[38] = 6'h35;
        mem[39] = 6'h28;
        mem[40] = 6'h16;
        mem[41] = 6'h07;
        mem[42] = 6'h05;
        mem[43] = 6'h3b;
        mem[44] = 6'h27;
        mem[45] = 6'h1f;
        mem[46] = 6'h3c;
        mem[47] = 6'h04;
        mem[48] = 6'h1b;
        mem[49] = 6'h02;
        mem[50] = 6'h17;
        mem[51] = 6'h0c;
        mem[52] = 6'h30;
        mem[53] = 6'h21;
        mem[54] = 6'h1c;
        mem[55] = 6'h2d;
        mem[56] = 6'h12;
        mem[57] = 6'h14;
        mem[58] = 6'h2e;
        mem[59] = 6'h18;
        mem[60] = 6'h36;
        mem[61] = 6'h31;
        mem[62] = 6'h0f;
        mem[63] = 6'h0e;
    end
endmodule

module odo_sbox_small2(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h13;
        mem[1] = 6'h3a;
        mem[2] = 6'h01;
        mem[3] = 6'h16;
        mem[4] = 6'h17;
        mem[5] = 6'h26;
        mem[6] = 6'h39;
        mem[7] = 6'h22;
        mem[8] = 6'h18;
        mem[9] = 6'h1c;
        mem[10] = 6'h3c;
        mem[11] = 6'h00;
        mem[12] = 6'h11;
        mem[13] = 6'h3e;
        mem[14] = 6'h12;
        mem[15] = 6'h14;
        mem[16] = 6'h30;
        mem[17] = 6'h1d;
        mem[18] = 6'h37;
        mem[19] = 6'h28;
        mem[20] = 6'h21;
        mem[21] = 6'h2a;
        mem[22] = 6'h19;
        mem[23] = 6'h0a;
        mem[24] = 6'h32;
        mem[25] = 6'h0b;
        mem[26] = 6'h1f;
        mem[27] = 6'h06;
        mem[28] = 6'h10;
        mem[29] = 6'h0c;
        mem[30] = 6'h38;
        mem[31] = 6'h2c;
        mem[32] = 6'h25;
        mem[33] = 6'h24;
        mem[34] = 6'h20;
        mem[35] = 6'h2e;
        mem[36] = 6'h3d;
        mem[37] = 6'h3b;
        mem[38] = 6'h33;
        mem[39] = 6'h0f;
        mem[40] = 6'h09;
        mem[41] = 6'h03;
        mem[42] = 6'h2d;
        mem[43] = 6'h1e;
        mem[44] = 6'h1a;
        mem[45] = 6'h3f;
        mem[46] = 6'h27;
        mem[47] = 6'h07;
        mem[48] = 6'h2b;
        mem[49] = 6'h04;
        mem[50] = 6'h36;
        mem[51] = 6'h0e;
        mem[52] = 6'h0d;
        mem[53] = 6'h15;
        mem[54] = 6'h05;
        mem[55] = 6'h02;
        mem[56] = 6'h29;
        mem[57] = 6'h1b;
        mem[58] = 6'h2f;
        mem[59] = 6'h23;
        mem[60] = 6'h08;
        mem[61] = 6'h34;
        mem[62] = 6'h31;
        mem[63] = 6'h35;
    end
endmodule

module odo_sbox_small3(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h38;
        mem[1] = 6'h3c;
        mem[2] = 6'h37;
        mem[3] = 6'h2b;
        mem[4] = 6'h05;
        mem[5] = 6'h14;
        mem[6] = 6'h09;
        mem[7] = 6'h1f;
        mem[8] = 6'h0e;
        mem[9] = 6'h12;
        mem[10] = 6'h35;
        mem[11] = 6'h0d;
        mem[12] = 6'h07;
        mem[13] = 6'h16;
        mem[14] = 6'h34;
        mem[15] = 6'h3d;
        mem[16] = 6'h10;
        mem[17] = 6'h29;
        mem[18] = 6'h31;
        mem[19] = 6'h28;
        mem[20] = 6'h24;
        mem[21] = 6'h13;
        mem[22] = 6'h11;
        mem[23] = 6'h1b;
        mem[24] = 6'h1e;
        mem[25] = 6'h21;
        mem[26] = 6'h22;
        mem[27] = 6'h3b;
        mem[28] = 6'h1a;
        mem[29] = 6'h30;
        mem[30] = 6'h0c;
        mem[31] = 6'h18;
        mem[32] = 6'h32;
        mem[33] = 6'h20;
        mem[34] = 6'h25;
        mem[35] = 6'h3f;
        mem[36] = 6'h06;
        mem[37] = 6'h03;
        mem[38] = 6'h3a;
        mem[39] = 6'h39;
        mem[40] = 6'h2a;
        mem[41] = 6'h27;
        mem[42] = 6'h23;
        mem[43] = 6'h2d;
        mem[44] = 6'h00;
        mem[45] = 6'h1d;
        mem[46] = 6'h3e;
        mem[47] = 6'h1c;
        mem[48] = 6'h2f;
        mem[49] = 6'h01;
        mem[50] = 6'h04;
        mem[51] = 6'h2e;
        mem[52] = 6'h2c;
        mem[53] = 6'h17;
        mem[54] = 6'h02;
        mem[55] = 6'h33;
        mem[56] = 6'h0f;
        mem[57] = 6'h19;
        mem[58] = 6'h0a;
        mem[59] = 6'h15;
        mem[60] = 6'h36;
        mem[61] = 6'h26;
        mem[62] = 6'h08;
        mem[63] = 6'h0b;
    end
endmodule

module odo_sbox_small4(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0a;
        mem[1] = 6'h39;
        mem[2] = 6'h15;
        mem[3] = 6'h03;
        mem[4] = 6'h1d;
        mem[5] = 6'h3d;
        mem[6] = 6'h00;
        mem[7] = 6'h34;
        mem[8] = 6'h06;
        mem[9] = 6'h25;
        mem[10] = 6'h0b;
        mem[11] = 6'h1f;
        mem[12] = 6'h26;
        mem[13] = 6'h0f;
        mem[14] = 6'h17;
        mem[15] = 6'h0d;
        mem[16] = 6'h05;
        mem[17] = 6'h0e;
        mem[18] = 6'h38;
        mem[19] = 6'h32;
        mem[20] = 6'h1a;
        mem[21] = 6'h33;
        mem[22] = 6'h31;
        mem[23] = 6'h07;
        mem[24] = 6'h1e;
        mem[25] = 6'h01;
        mem[26] = 6'h19;
        mem[27] = 6'h2f;
        mem[28] = 6'h2a;
        mem[29] = 6'h2b;
        mem[30] = 6'h11;
        mem[31] = 6'h29;
        mem[32] = 6'h08;
        mem[33] = 6'h10;
        mem[34] = 6'h22;
        mem[35] = 6'h21;
        mem[36] = 6'h12;
        mem[37] = 6'h36;
        mem[38] = 6'h02;
        mem[39] = 6'h3c;
        mem[40] = 6'h04;
        mem[41] = 6'h28;
        mem[42] = 6'h3f;
        mem[43] = 6'h35;
        mem[44] = 6'h3a;
        mem[45] = 6'h2e;
        mem[46] = 6'h37;
        mem[47] = 6'h2d;
        mem[48] = 6'h1c;
        mem[49] = 6'h2c;
        mem[50] = 6'h23;
        mem[51] = 6'h1b;
        mem[52] = 6'h16;
        mem[53] = 6'h3b;
        mem[54] = 6'h24;
        mem[55] = 6'h13;
        mem[56] = 6'h18;
        mem[57] = 6'h0c;
        mem[58] = 6'h3e;
        mem[59] = 6'h20;
        mem[60] = 6'h14;
        mem[61] = 6'h09;
        mem[62] = 6'h30;
        mem[63] = 6'h27;
    end
endmodule

module odo_sbox_small5(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h31;
        mem[1] = 6'h2e;
        mem[2] = 6'h09;
        mem[3] = 6'h08;
        mem[4] = 6'h2a;
        mem[5] = 6'h04;
        mem[6] = 6'h29;
        mem[7] = 6'h25;
        mem[8] = 6'h1d;
        mem[9] = 6'h24;
        mem[10] = 6'h01;
        mem[11] = 6'h10;
        mem[12] = 6'h0b;
        mem[13] = 6'h1e;
        mem[14] = 6'h03;
        mem[15] = 6'h07;
        mem[16] = 6'h38;
        mem[17] = 6'h1a;
        mem[18] = 6'h02;
        mem[19] = 6'h3d;
        mem[20] = 6'h3b;
        mem[21] = 6'h15;
        mem[22] = 6'h1c;
        mem[23] = 6'h0e;
        mem[24] = 6'h2f;
        mem[25] = 6'h18;
        mem[26] = 6'h39;
        mem[27] = 6'h1f;
        mem[28] = 6'h33;
        mem[29] = 6'h34;
        mem[30] = 6'h32;
        mem[31] = 6'h0f;
        mem[32] = 6'h14;
        mem[33] = 6'h05;
        mem[34] = 6'h1b;
        mem[35] = 6'h23;
        mem[36] = 6'h06;
        mem[37] = 6'h2b;
        mem[38] = 6'h0c;
        mem[39] = 6'h19;
        mem[40] = 6'h0a;
        mem[41] = 6'h37;
        mem[42] = 6'h30;
        mem[43] = 6'h28;
        mem[44] = 6'h2d;
        mem[45] = 6'h17;
        mem[46] = 6'h35;
        mem[47] = 6'h26;
        mem[48] = 6'h3a;
        mem[49] = 6'h20;
        mem[50] = 6'h11;
        mem[51] = 6'h12;
        mem[52] = 6'h3f;
        mem[53] = 6'h00;
        mem[54] = 6'h27;
        mem[55] = 6'h2c;
        mem[56] = 6'h22;
        mem[57] = 6'h3e;
        mem[58] = 6'h0d;
        mem[59] = 6'h16;
        mem[60] = 6'h3c;
        mem[61] = 6'h36;
        mem[62] = 6'h21;
        mem[63] = 6'h13;
    end
endmodule

module odo_sbox_small6(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h35;
        mem[1] = 6'h04;
        mem[2] = 6'h0f;
        mem[3] = 6'h31;
        mem[4] = 6'h32;
        mem[5] = 6'h03;
        mem[6] = 6'h1a;
        mem[7] = 6'h01;
        mem[8] = 6'h16;
        mem[9] = 6'h26;
        mem[10] = 6'h2a;
        mem[11] = 6'h29;
        mem[12] = 6'h27;
        mem[13] = 6'h13;
        mem[14] = 6'h12;
        mem[15] = 6'h3c;
        mem[16] = 6'h1d;
        mem[17] = 6'h3d;
        mem[18] = 6'h36;
        mem[19] = 6'h34;
        mem[20] = 6'h06;
        mem[21] = 6'h37;
        mem[22] = 6'h28;
        mem[23] = 6'h2b;
        mem[24] = 6'h3a;
        mem[25] = 6'h0d;
        mem[26] = 6'h1c;
        mem[27] = 6'h02;
        mem[28] = 6'h00;
        mem[29] = 6'h33;
        mem[30] = 6'h0c;
        mem[31] = 6'h3b;
        mem[32] = 6'h24;
        mem[33] = 6'h3f;
        mem[34] = 6'h2f;
        mem[35] = 6'h1e;
        mem[36] = 6'h2e;
        mem[37] = 6'h2d;
        mem[38] = 6'h0a;
        mem[39] = 6'h17;
        mem[40] = 6'h20;
        mem[41] = 6'h0b;
        mem[42] = 6'h15;
        mem[43] = 6'h1f;
        mem[44] = 6'h14;
        mem[45] = 6'h3e;
        mem[46] = 6'h25;
        mem[47] = 6'h11;
        mem[48] = 6'h38;
        mem[49] = 6'h09;
        mem[50] = 6'h23;
        mem[51] = 6'h0e;
        mem[52] = 6'h1b;
        mem[53] = 6'h18;
        mem[54] = 6'h08;
        mem[55] = 6'h19;
        mem[56] = 6'h2c;
        mem[57] = 6'h05;
        mem[58] = 6'h21;
        mem[59] = 6'h39;
        mem[60] = 6'h07;
        mem[61] = 6'h10;
        mem[62] = 6'h30;
        mem[63] = 6'h22;
    end
endmodule

module odo_sbox_small7(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h22;
        mem[1] = 6'h26;
        mem[2] = 6'h19;
        mem[3] = 6'h20;
        mem[4] = 6'h3e;
        mem[5] = 6'h2a;
        mem[6] = 6'h1b;
        mem[7] = 6'h0f;
        mem[8] = 6'h14;
        mem[9] = 6'h11;
        mem[10] = 6'h1d;
        mem[11] = 6'h33;
        mem[12] = 6'h00;
        mem[13] = 6'h29;
        mem[14] = 6'h1c;
        mem[15] = 6'h35;
        mem[16] = 6'h04;
        mem[17] = 6'h2d;
        mem[18] = 6'h1a;
        mem[19] = 6'h32;
        mem[20] = 6'h38;
        mem[21] = 6'h13;
        mem[22] = 6'h37;
        mem[23] = 6'h2c;
        mem[24] = 6'h3a;
        mem[25] = 6'h09;
        mem[26] = 6'h0a;
        mem[27] = 6'h03;
        mem[28] = 6'h01;
        mem[29] = 6'h1e;
        mem[30] = 6'h16;
        mem[31] = 6'h3b;
        mem[32] = 6'h2b;
        mem[33] = 6'h08;
        mem[34] = 6'h3c;
        mem[35] = 6'h0c;
        mem[36] = 6'h1f;
        mem[37] = 6'h2f;
        mem[38] = 6'h27;
        mem[39] = 6'h12;
        mem[40] = 6'h2e;
        mem[41] = 6'h23;
        mem[42] = 6'h3f;
        mem[43] = 6'h0b;
        mem[44] = 6'h0e;
        mem[45] = 6'h24;
        mem[46] = 6'h39;
        mem[47] = 6'h06;
        mem[48] = 6'h25;
        mem[49] = 6'h31;
        mem[50] = 6'h02;
        mem[51] = 6'h30;
        mem[52] = 6'h17;
        mem[53] = 6'h28;
        mem[54] = 6'h36;
        mem[55] = 6'h21;
        mem[56] = 6'h0d;
        mem[57] = 6'h15;
        mem[58] = 6'h10;
        mem[59] = 6'h07;
        mem[60] = 6'h34;
        mem[61] = 6'h05;
        mem[62] = 6'h18;
        mem[63] = 6'h3d;
    end
endmodule

module odo_sbox_small8(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h06;
        mem[1] = 6'h2e;
        mem[2] = 6'h19;
        mem[3] = 6'h24;
        mem[4] = 6'h31;
        mem[5] = 6'h20;
        mem[6] = 6'h0a;
        mem[7] = 6'h2a;
        mem[8] = 6'h3c;
        mem[9] = 6'h09;
        mem[10] = 6'h2b;
        mem[11] = 6'h34;
        mem[12] = 6'h37;
        mem[13] = 6'h0b;
        mem[14] = 6'h1c;
        mem[15] = 6'h3b;
        mem[16] = 6'h21;
        mem[17] = 6'h04;
        mem[18] = 6'h3d;
        mem[19] = 6'h0c;
        mem[20] = 6'h28;
        mem[21] = 6'h1a;
        mem[22] = 6'h18;
        mem[23] = 6'h15;
        mem[24] = 6'h05;
        mem[25] = 6'h1d;
        mem[26] = 6'h0f;
        mem[27] = 6'h00;
        mem[28] = 6'h02;
        mem[29] = 6'h2f;
        mem[30] = 6'h13;
        mem[31] = 6'h2d;
        mem[32] = 6'h30;
        mem[33] = 6'h1e;
        mem[34] = 6'h2c;
        mem[35] = 6'h0e;
        mem[36] = 6'h36;
        mem[37] = 6'h1b;
        mem[38] = 6'h27;
        mem[39] = 6'h03;
        mem[40] = 6'h3e;
        mem[41] = 6'h35;
        mem[42] = 6'h17;
        mem[43] = 6'h38;
        mem[44] = 6'h16;
        mem[45] = 6'h33;
        mem[46] = 6'h12;
        mem[47] = 6'h29;
        mem[48] = 6'h39;
        mem[49] = 6'h08;
        mem[50] = 6'h3f;
        mem[51] = 6'h0d;
        mem[52] = 6'h11;
        mem[53] = 6'h07;
        mem[54] = 6'h10;
        mem[55] = 6'h01;
        mem[56] = 6'h23;
        mem[57] = 6'h1f;
        mem[58] = 6'h26;
        mem[59] = 6'h14;
        mem[60] = 6'h32;
        mem[61] = 6'h3a;
        mem[62] = 6'h22;
        mem[63] = 6'h25;
    end
endmodule

module odo_sbox_small9(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1a;
        mem[1] = 6'h15;
        mem[2] = 6'h06;
        mem[3] = 6'h11;
        mem[4] = 6'h2b;
        mem[5] = 6'h0d;
        mem[6] = 6'h1b;
        mem[7] = 6'h00;
        mem[8] = 6'h27;
        mem[9] = 6'h28;
        mem[10] = 6'h3e;
        mem[11] = 6'h25;
        mem[12] = 6'h32;
        mem[13] = 6'h2d;
        mem[14] = 6'h30;
        mem[15] = 6'h22;
        mem[16] = 6'h13;
        mem[17] = 6'h26;
        mem[18] = 6'h02;
        mem[19] = 6'h12;
        mem[20] = 6'h01;
        mem[21] = 6'h1f;
        mem[22] = 6'h16;
        mem[23] = 6'h0a;
        mem[24] = 6'h14;
        mem[25] = 6'h23;
        mem[26] = 6'h3f;
        mem[27] = 6'h20;
        mem[28] = 6'h29;
        mem[29] = 6'h0c;
        mem[30] = 6'h38;
        mem[31] = 6'h36;
        mem[32] = 6'h34;
        mem[33] = 6'h19;
        mem[34] = 6'h31;
        mem[35] = 6'h3a;
        mem[36] = 6'h09;
        mem[37] = 6'h0b;
        mem[38] = 6'h05;
        mem[39] = 6'h1e;
        mem[40] = 6'h1d;
        mem[41] = 6'h0e;
        mem[42] = 6'h39;
        mem[43] = 6'h35;
        mem[44] = 6'h18;
        mem[45] = 6'h10;
        mem[46] = 6'h03;
        mem[47] = 6'h07;
        mem[48] = 6'h17;
        mem[49] = 6'h37;
        mem[50] = 6'h0f;
        mem[51] = 6'h1c;
        mem[52] = 6'h2a;
        mem[53] = 6'h3c;
        mem[54] = 6'h3b;
        mem[55] = 6'h33;
        mem[56] = 6'h2e;
        mem[57] = 6'h2f;
        mem[58] = 6'h2c;
        mem[59] = 6'h08;
        mem[60] = 6'h21;
        mem[61] = 6'h3d;
        mem[62] = 6'h04;
        mem[63] = 6'h24;
    end
endmodule

module odo_sbox_small10(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1e;
        mem[1] = 6'h18;
        mem[2] = 6'h20;
        mem[3] = 6'h19;
        mem[4] = 6'h28;
        mem[5] = 6'h3e;
        mem[6] = 6'h36;
        mem[7] = 6'h2a;
        mem[8] = 6'h29;
        mem[9] = 6'h10;
        mem[10] = 6'h01;
        mem[11] = 6'h39;
        mem[12] = 6'h05;
        mem[13] = 6'h35;
        mem[14] = 6'h15;
        mem[15] = 6'h1c;
        mem[16] = 6'h00;
        mem[17] = 6'h06;
        mem[18] = 6'h14;
        mem[19] = 6'h09;
        mem[20] = 6'h17;
        mem[21] = 6'h3d;
        mem[22] = 6'h13;
        mem[23] = 6'h0d;
        mem[24] = 6'h08;
        mem[25] = 6'h3c;
        mem[26] = 6'h26;
        mem[27] = 6'h16;
        mem[28] = 6'h12;
        mem[29] = 6'h2b;
        mem[30] = 6'h0b;
        mem[31] = 6'h38;
        mem[32] = 6'h23;
        mem[33] = 6'h2e;
        mem[34] = 6'h1a;
        mem[35] = 6'h0c;
        mem[36] = 6'h3f;
        mem[37] = 6'h1d;
        mem[38] = 6'h30;
        mem[39] = 6'h02;
        mem[40] = 6'h24;
        mem[41] = 6'h33;
        mem[42] = 6'h0e;
        mem[43] = 6'h11;
        mem[44] = 6'h0a;
        mem[45] = 6'h1b;
        mem[46] = 6'h2f;
        mem[47] = 6'h2d;
        mem[48] = 6'h27;
        mem[49] = 6'h31;
        mem[50] = 6'h37;
        mem[51] = 6'h22;
        mem[52] = 6'h34;
        mem[53] = 6'h07;
        mem[54] = 6'h3b;
        mem[55] = 6'h04;
        mem[56] = 6'h32;
        mem[57] = 6'h2c;
        mem[58] = 6'h25;
        mem[59] = 6'h1f;
        mem[60] = 6'h21;
        mem[61] = 6'h03;
        mem[62] = 6'h0f;
        mem[63] = 6'h3a;
    end
endmodule

module odo_sbox_small11(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h35;
        mem[1] = 6'h04;
        mem[2] = 6'h32;
        mem[3] = 6'h38;
        mem[4] = 6'h06;
        mem[5] = 6'h0b;
        mem[6] = 6'h31;
        mem[7] = 6'h2e;
        mem[8] = 6'h30;
        mem[9] = 6'h20;
        mem[10] = 6'h03;
        mem[11] = 6'h1c;
        mem[12] = 6'h00;
        mem[13] = 6'h1b;
        mem[14] = 6'h25;
        mem[15] = 6'h33;
        mem[16] = 6'h0a;
        mem[17] = 6'h02;
        mem[18] = 6'h37;
        mem[19] = 6'h3a;
        mem[20] = 6'h2d;
        mem[21] = 6'h0d;
        mem[22] = 6'h11;
        mem[23] = 6'h29;
        mem[24] = 6'h26;
        mem[25] = 6'h3e;
        mem[26] = 6'h2f;
        mem[27] = 6'h3d;
        mem[28] = 6'h13;
        mem[29] = 6'h0c;
        mem[30] = 6'h0e;
        mem[31] = 6'h24;
        mem[32] = 6'h21;
        mem[33] = 6'h2a;
        mem[34] = 6'h22;
        mem[35] = 6'h36;
        mem[36] = 6'h1e;
        mem[37] = 6'h1d;
        mem[38] = 6'h16;
        mem[39] = 6'h1f;
        mem[40] = 6'h01;
        mem[41] = 6'h3b;
        mem[42] = 6'h09;
        mem[43] = 6'h27;
        mem[44] = 6'h08;
        mem[45] = 6'h2c;
        mem[46] = 6'h05;
        mem[47] = 6'h28;
        mem[48] = 6'h18;
        mem[49] = 6'h2b;
        mem[50] = 6'h23;
        mem[51] = 6'h1a;
        mem[52] = 6'h12;
        mem[53] = 6'h39;
        mem[54] = 6'h10;
        mem[55] = 6'h14;
        mem[56] = 6'h17;
        mem[57] = 6'h3f;
        mem[58] = 6'h34;
        mem[59] = 6'h07;
        mem[60] = 6'h15;
        mem[61] = 6'h3c;
        mem[62] = 6'h0f;
        mem[63] = 6'h19;
    end
endmodule

module odo_sbox_small12(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2c;
        mem[1] = 6'h04;
        mem[2] = 6'h24;
        mem[3] = 6'h05;
        mem[4] = 6'h2a;
        mem[5] = 6'h37;
        mem[6] = 6'h07;
        mem[7] = 6'h38;
        mem[8] = 6'h3f;
        mem[9] = 6'h0e;
        mem[10] = 6'h1e;
        mem[11] = 6'h21;
        mem[12] = 6'h32;
        mem[13] = 6'h1a;
        mem[14] = 6'h0c;
        mem[15] = 6'h35;
        mem[16] = 6'h36;
        mem[17] = 6'h26;
        mem[18] = 6'h30;
        mem[19] = 6'h02;
        mem[20] = 6'h0a;
        mem[21] = 6'h00;
        mem[22] = 6'h12;
        mem[23] = 6'h29;
        mem[24] = 6'h03;
        mem[25] = 6'h10;
        mem[26] = 6'h0b;
        mem[27] = 6'h0d;
        mem[28] = 6'h14;
        mem[29] = 6'h09;
        mem[30] = 6'h17;
        mem[31] = 6'h19;
        mem[32] = 6'h20;
        mem[33] = 6'h39;
        mem[34] = 6'h25;
        mem[35] = 6'h33;
        mem[36] = 6'h3e;
        mem[37] = 6'h0f;
        mem[38] = 6'h11;
        mem[39] = 6'h34;
        mem[40] = 6'h16;
        mem[41] = 6'h1d;
        mem[42] = 6'h27;
        mem[43] = 6'h2f;
        mem[44] = 6'h3b;
        mem[45] = 6'h18;
        mem[46] = 6'h2e;
        mem[47] = 6'h08;
        mem[48] = 6'h2b;
        mem[49] = 6'h06;
        mem[50] = 6'h15;
        mem[51] = 6'h2d;
        mem[52] = 6'h01;
        mem[53] = 6'h1f;
        mem[54] = 6'h3a;
        mem[55] = 6'h28;
        mem[56] = 6'h3c;
        mem[57] = 6'h13;
        mem[58] = 6'h22;
        mem[59] = 6'h1b;
        mem[60] = 6'h31;
        mem[61] = 6'h3d;
        mem[62] = 6'h23;
        mem[63] = 6'h1c;
    end
endmodule

module odo_sbox_small13(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0c;
        mem[1] = 6'h28;
        mem[2] = 6'h17;
        mem[3] = 6'h29;
        mem[4] = 6'h37;
        mem[5] = 6'h20;
        mem[6] = 6'h1b;
        mem[7] = 6'h3a;
        mem[8] = 6'h03;
        mem[9] = 6'h19;
        mem[10] = 6'h0f;
        mem[11] = 6'h0b;
        mem[12] = 6'h09;
        mem[13] = 6'h1d;
        mem[14] = 6'h30;
        mem[15] = 6'h35;
        mem[16] = 6'h27;
        mem[17] = 6'h12;
        mem[18] = 6'h1f;
        mem[19] = 6'h33;
        mem[20] = 6'h2a;
        mem[21] = 6'h21;
        mem[22] = 6'h08;
        mem[23] = 6'h11;
        mem[24] = 6'h3e;
        mem[25] = 6'h1a;
        mem[26] = 6'h2d;
        mem[27] = 6'h06;
        mem[28] = 6'h31;
        mem[29] = 6'h3c;
        mem[30] = 6'h39;
        mem[31] = 6'h2b;
        mem[32] = 6'h34;
        mem[33] = 6'h0e;
        mem[34] = 6'h38;
        mem[35] = 6'h3b;
        mem[36] = 6'h05;
        mem[37] = 6'h15;
        mem[38] = 6'h16;
        mem[39] = 6'h0a;
        mem[40] = 6'h23;
        mem[41] = 6'h24;
        mem[42] = 6'h14;
        mem[43] = 6'h2c;
        mem[44] = 6'h2e;
        mem[45] = 6'h1e;
        mem[46] = 6'h26;
        mem[47] = 6'h00;
        mem[48] = 6'h36;
        mem[49] = 6'h13;
        mem[50] = 6'h01;
        mem[51] = 6'h1c;
        mem[52] = 6'h3f;
        mem[53] = 6'h04;
        mem[54] = 6'h10;
        mem[55] = 6'h25;
        mem[56] = 6'h18;
        mem[57] = 6'h3d;
        mem[58] = 6'h22;
        mem[59] = 6'h0d;
        mem[60] = 6'h2f;
        mem[61] = 6'h02;
        mem[62] = 6'h07;
        mem[63] = 6'h32;
    end
endmodule

module odo_sbox_small14(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1a;
        mem[1] = 6'h2a;
        mem[2] = 6'h10;
        mem[3] = 6'h09;
        mem[4] = 6'h30;
        mem[5] = 6'h1f;
        mem[6] = 6'h11;
        mem[7] = 6'h31;
        mem[8] = 6'h16;
        mem[9] = 6'h33;
        mem[10] = 6'h14;
        mem[11] = 6'h3c;
        mem[12] = 6'h1d;
        mem[13] = 6'h35;
        mem[14] = 6'h19;
        mem[15] = 6'h17;
        mem[16] = 6'h04;
        mem[17] = 6'h02;
        mem[18] = 6'h03;
        mem[19] = 6'h26;
        mem[20] = 6'h24;
        mem[21] = 6'h3f;
        mem[22] = 6'h0f;
        mem[23] = 6'h1e;
        mem[24] = 6'h36;
        mem[25] = 6'h0e;
        mem[26] = 6'h21;
        mem[27] = 6'h08;
        mem[28] = 6'h27;
        mem[29] = 6'h20;
        mem[30] = 6'h2e;
        mem[31] = 6'h0a;
        mem[32] = 6'h06;
        mem[33] = 6'h23;
        mem[34] = 6'h34;
        mem[35] = 6'h07;
        mem[36] = 6'h1b;
        mem[37] = 6'h0b;
        mem[38] = 6'h2d;
        mem[39] = 6'h37;
        mem[40] = 6'h29;
        mem[41] = 6'h25;
        mem[42] = 6'h2c;
        mem[43] = 6'h3b;
        mem[44] = 6'h0d;
        mem[45] = 6'h2b;
        mem[46] = 6'h05;
        mem[47] = 6'h3a;
        mem[48] = 6'h32;
        mem[49] = 6'h3e;
        mem[50] = 6'h00;
        mem[51] = 6'h39;
        mem[52] = 6'h38;
        mem[53] = 6'h01;
        mem[54] = 6'h1c;
        mem[55] = 6'h22;
        mem[56] = 6'h2f;
        mem[57] = 6'h13;
        mem[58] = 6'h15;
        mem[59] = 6'h0c;
        mem[60] = 6'h3d;
        mem[61] = 6'h28;
        mem[62] = 6'h18;
        mem[63] = 6'h12;
    end
endmodule

module odo_sbox_small15(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h18;
        mem[1] = 6'h11;
        mem[2] = 6'h1d;
        mem[3] = 6'h1c;
        mem[4] = 6'h23;
        mem[5] = 6'h3d;
        mem[6] = 6'h15;
        mem[7] = 6'h34;
        mem[8] = 6'h20;
        mem[9] = 6'h0e;
        mem[10] = 6'h16;
        mem[11] = 6'h02;
        mem[12] = 6'h3b;
        mem[13] = 6'h04;
        mem[14] = 6'h19;
        mem[15] = 6'h36;
        mem[16] = 6'h25;
        mem[17] = 6'h0b;
        mem[18] = 6'h3f;
        mem[19] = 6'h0f;
        mem[20] = 6'h2d;
        mem[21] = 6'h29;
        mem[22] = 6'h07;
        mem[23] = 6'h13;
        mem[24] = 6'h14;
        mem[25] = 6'h39;
        mem[26] = 6'h10;
        mem[27] = 6'h24;
        mem[28] = 6'h3e;
        mem[29] = 6'h22;
        mem[30] = 6'h0d;
        mem[31] = 6'h2c;
        mem[32] = 6'h00;
        mem[33] = 6'h33;
        mem[34] = 6'h26;
        mem[35] = 6'h01;
        mem[36] = 6'h1a;
        mem[37] = 6'h1b;
        mem[38] = 6'h3c;
        mem[39] = 6'h17;
        mem[40] = 6'h09;
        mem[41] = 6'h1f;
        mem[42] = 6'h2f;
        mem[43] = 6'h2e;
        mem[44] = 6'h2a;
        mem[45] = 6'h28;
        mem[46] = 6'h32;
        mem[47] = 6'h0a;
        mem[48] = 6'h3a;
        mem[49] = 6'h38;
        mem[50] = 6'h21;
        mem[51] = 6'h2b;
        mem[52] = 6'h27;
        mem[53] = 6'h31;
        mem[54] = 6'h0c;
        mem[55] = 6'h35;
        mem[56] = 6'h12;
        mem[57] = 6'h37;
        mem[58] = 6'h30;
        mem[59] = 6'h08;
        mem[60] = 6'h06;
        mem[61] = 6'h05;
        mem[62] = 6'h03;
        mem[63] = 6'h1e;
    end
endmodule

module odo_sbox_small16(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3a;
        mem[1] = 6'h31;
        mem[2] = 6'h02;
        mem[3] = 6'h17;
        mem[4] = 6'h29;
        mem[5] = 6'h3f;
        mem[6] = 6'h2d;
        mem[7] = 6'h23;
        mem[8] = 6'h2a;
        mem[9] = 6'h0a;
        mem[10] = 6'h1e;
        mem[11] = 6'h1d;
        mem[12] = 6'h2c;
        mem[13] = 6'h2e;
        mem[14] = 6'h3e;
        mem[15] = 6'h34;
        mem[16] = 6'h20;
        mem[17] = 6'h25;
        mem[18] = 6'h2b;
        mem[19] = 6'h03;
        mem[20] = 6'h3d;
        mem[21] = 6'h10;
        mem[22] = 6'h16;
        mem[23] = 6'h01;
        mem[24] = 6'h08;
        mem[25] = 6'h28;
        mem[26] = 6'h3c;
        mem[27] = 6'h12;
        mem[28] = 6'h13;
        mem[29] = 6'h36;
        mem[30] = 6'h00;
        mem[31] = 6'h26;
        mem[32] = 6'h22;
        mem[33] = 6'h14;
        mem[34] = 6'h1b;
        mem[35] = 6'h09;
        mem[36] = 6'h32;
        mem[37] = 6'h0f;
        mem[38] = 6'h0e;
        mem[39] = 6'h38;
        mem[40] = 6'h0d;
        mem[41] = 6'h0b;
        mem[42] = 6'h27;
        mem[43] = 6'h33;
        mem[44] = 6'h07;
        mem[45] = 6'h1c;
        mem[46] = 6'h11;
        mem[47] = 6'h05;
        mem[48] = 6'h30;
        mem[49] = 6'h21;
        mem[50] = 6'h1f;
        mem[51] = 6'h3b;
        mem[52] = 6'h19;
        mem[53] = 6'h24;
        mem[54] = 6'h2f;
        mem[55] = 6'h39;
        mem[56] = 6'h15;
        mem[57] = 6'h0c;
        mem[58] = 6'h06;
        mem[59] = 6'h18;
        mem[60] = 6'h35;
        mem[61] = 6'h37;
        mem[62] = 6'h1a;
        mem[63] = 6'h04;
    end
endmodule

module odo_sbox_small17(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h02;
        mem[1] = 6'h09;
        mem[2] = 6'h17;
        mem[3] = 6'h04;
        mem[4] = 6'h3e;
        mem[5] = 6'h15;
        mem[6] = 6'h05;
        mem[7] = 6'h1c;
        mem[8] = 6'h20;
        mem[9] = 6'h3f;
        mem[10] = 6'h00;
        mem[11] = 6'h1f;
        mem[12] = 6'h37;
        mem[13] = 6'h3c;
        mem[14] = 6'h0f;
        mem[15] = 6'h25;
        mem[16] = 6'h32;
        mem[17] = 6'h39;
        mem[18] = 6'h19;
        mem[19] = 6'h1b;
        mem[20] = 6'h26;
        mem[21] = 6'h1d;
        mem[22] = 6'h34;
        mem[23] = 6'h2c;
        mem[24] = 6'h0e;
        mem[25] = 6'h1a;
        mem[26] = 6'h06;
        mem[27] = 6'h35;
        mem[28] = 6'h36;
        mem[29] = 6'h38;
        mem[30] = 6'h12;
        mem[31] = 6'h33;
        mem[32] = 6'h0c;
        mem[33] = 6'h2a;
        mem[34] = 6'h21;
        mem[35] = 6'h24;
        mem[36] = 6'h0d;
        mem[37] = 6'h03;
        mem[38] = 6'h2d;
        mem[39] = 6'h01;
        mem[40] = 6'h13;
        mem[41] = 6'h0b;
        mem[42] = 6'h22;
        mem[43] = 6'h10;
        mem[44] = 6'h3b;
        mem[45] = 6'h27;
        mem[46] = 6'h3a;
        mem[47] = 6'h3d;
        mem[48] = 6'h23;
        mem[49] = 6'h30;
        mem[50] = 6'h31;
        mem[51] = 6'h18;
        mem[52] = 6'h1e;
        mem[53] = 6'h2b;
        mem[54] = 6'h11;
        mem[55] = 6'h14;
        mem[56] = 6'h2f;
        mem[57] = 6'h08;
        mem[58] = 6'h28;
        mem[59] = 6'h2e;
        mem[60] = 6'h29;
        mem[61] = 6'h0a;
        mem[62] = 6'h07;
        mem[63] = 6'h16;
    end
endmodule

module odo_sbox_small18(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h05;
        mem[1] = 6'h27;
        mem[2] = 6'h2f;
        mem[3] = 6'h30;
        mem[4] = 6'h25;
        mem[5] = 6'h24;
        mem[6] = 6'h02;
        mem[7] = 6'h1e;
        mem[8] = 6'h1b;
        mem[9] = 6'h33;
        mem[10] = 6'h1f;
        mem[11] = 6'h3e;
        mem[12] = 6'h21;
        mem[13] = 6'h01;
        mem[14] = 6'h11;
        mem[15] = 6'h17;
        mem[16] = 6'h3a;
        mem[17] = 6'h07;
        mem[18] = 6'h1c;
        mem[19] = 6'h15;
        mem[20] = 6'h31;
        mem[21] = 6'h38;
        mem[22] = 6'h06;
        mem[23] = 6'h29;
        mem[24] = 6'h37;
        mem[25] = 6'h2a;
        mem[26] = 6'h35;
        mem[27] = 6'h2c;
        mem[28] = 6'h20;
        mem[29] = 6'h10;
        mem[30] = 6'h22;
        mem[31] = 6'h0b;
        mem[32] = 6'h12;
        mem[33] = 6'h36;
        mem[34] = 6'h1a;
        mem[35] = 6'h23;
        mem[36] = 6'h1d;
        mem[37] = 6'h39;
        mem[38] = 6'h19;
        mem[39] = 6'h34;
        mem[40] = 6'h2b;
        mem[41] = 6'h0f;
        mem[42] = 6'h3f;
        mem[43] = 6'h14;
        mem[44] = 6'h3d;
        mem[45] = 6'h0e;
        mem[46] = 6'h0a;
        mem[47] = 6'h0d;
        mem[48] = 6'h32;
        mem[49] = 6'h28;
        mem[50] = 6'h13;
        mem[51] = 6'h03;
        mem[52] = 6'h09;
        mem[53] = 6'h26;
        mem[54] = 6'h3c;
        mem[55] = 6'h00;
        mem[56] = 6'h0c;
        mem[57] = 6'h2d;
        mem[58] = 6'h16;
        mem[59] = 6'h04;
        mem[60] = 6'h08;
        mem[61] = 6'h18;
        mem[62] = 6'h3b;
        mem[63] = 6'h2e;
    end
endmodule

module odo_sbox_small19(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h05;
        mem[1] = 6'h3d;
        mem[2] = 6'h1c;
        mem[3] = 6'h26;
        mem[4] = 6'h1e;
        mem[5] = 6'h13;
        mem[6] = 6'h0b;
        mem[7] = 6'h02;
        mem[8] = 6'h03;
        mem[9] = 6'h10;
        mem[10] = 6'h2a;
        mem[11] = 6'h0d;
        mem[12] = 6'h2d;
        mem[13] = 6'h24;
        mem[14] = 6'h34;
        mem[15] = 6'h18;
        mem[16] = 6'h1f;
        mem[17] = 6'h3a;
        mem[18] = 6'h19;
        mem[19] = 6'h04;
        mem[20] = 6'h1a;
        mem[21] = 6'h01;
        mem[22] = 6'h2f;
        mem[23] = 6'h3f;
        mem[24] = 6'h0c;
        mem[25] = 6'h39;
        mem[26] = 6'h0a;
        mem[27] = 6'h37;
        mem[28] = 6'h06;
        mem[29] = 6'h15;
        mem[30] = 6'h07;
        mem[31] = 6'h36;
        mem[32] = 6'h33;
        mem[33] = 6'h11;
        mem[34] = 6'h00;
        mem[35] = 6'h32;
        mem[36] = 6'h3c;
        mem[37] = 6'h2e;
        mem[38] = 6'h0f;
        mem[39] = 6'h21;
        mem[40] = 6'h2b;
        mem[41] = 6'h1d;
        mem[42] = 6'h25;
        mem[43] = 6'h09;
        mem[44] = 6'h22;
        mem[45] = 6'h31;
        mem[46] = 6'h38;
        mem[47] = 6'h23;
        mem[48] = 6'h2c;
        mem[49] = 6'h27;
        mem[50] = 6'h16;
        mem[51] = 6'h30;
        mem[52] = 6'h17;
        mem[53] = 6'h14;
        mem[54] = 6'h0e;
        mem[55] = 6'h29;
        mem[56] = 6'h20;
        mem[57] = 6'h12;
        mem[58] = 6'h3b;
        mem[59] = 6'h08;
        mem[60] = 6'h35;
        mem[61] = 6'h3e;
        mem[62] = 6'h28;
        mem[63] = 6'h1b;
    end
endmodule

module odo_sbox_small20(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h05;
        mem[1] = 6'h12;
        mem[2] = 6'h23;
        mem[3] = 6'h2a;
        mem[4] = 6'h14;
        mem[5] = 6'h2d;
        mem[6] = 6'h31;
        mem[7] = 6'h1b;
        mem[8] = 6'h01;
        mem[9] = 6'h21;
        mem[10] = 6'h35;
        mem[11] = 6'h19;
        mem[12] = 6'h2b;
        mem[13] = 6'h09;
        mem[14] = 6'h11;
        mem[15] = 6'h29;
        mem[16] = 6'h0f;
        mem[17] = 6'h25;
        mem[18] = 6'h02;
        mem[19] = 6'h39;
        mem[20] = 6'h3e;
        mem[21] = 6'h08;
        mem[22] = 6'h38;
        mem[23] = 6'h0e;
        mem[24] = 6'h0b;
        mem[25] = 6'h37;
        mem[26] = 6'h30;
        mem[27] = 6'h34;
        mem[28] = 6'h10;
        mem[29] = 6'h07;
        mem[30] = 6'h32;
        mem[31] = 6'h0c;
        mem[32] = 6'h24;
        mem[33] = 6'h20;
        mem[34] = 6'h36;
        mem[35] = 6'h16;
        mem[36] = 6'h3b;
        mem[37] = 6'h06;
        mem[38] = 6'h00;
        mem[39] = 6'h13;
        mem[40] = 6'h1e;
        mem[41] = 6'h1a;
        mem[42] = 6'h0d;
        mem[43] = 6'h3c;
        mem[44] = 6'h2e;
        mem[45] = 6'h28;
        mem[46] = 6'h0a;
        mem[47] = 6'h1f;
        mem[48] = 6'h04;
        mem[49] = 6'h3f;
        mem[50] = 6'h3d;
        mem[51] = 6'h3a;
        mem[52] = 6'h1c;
        mem[53] = 6'h1d;
        mem[54] = 6'h33;
        mem[55] = 6'h17;
        mem[56] = 6'h15;
        mem[57] = 6'h18;
        mem[58] = 6'h26;
        mem[59] = 6'h2c;
        mem[60] = 6'h27;
        mem[61] = 6'h2f;
        mem[62] = 6'h03;
        mem[63] = 6'h22;
    end
endmodule

module odo_sbox_small21(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h22;
        mem[1] = 6'h25;
        mem[2] = 6'h04;
        mem[3] = 6'h10;
        mem[4] = 6'h38;
        mem[5] = 6'h03;
        mem[6] = 6'h1e;
        mem[7] = 6'h1b;
        mem[8] = 6'h0d;
        mem[9] = 6'h3b;
        mem[10] = 6'h1d;
        mem[11] = 6'h34;
        mem[12] = 6'h2a;
        mem[13] = 6'h28;
        mem[14] = 6'h29;
        mem[15] = 6'h3c;
        mem[16] = 6'h14;
        mem[17] = 6'h0f;
        mem[18] = 6'h39;
        mem[19] = 6'h30;
        mem[20] = 6'h1f;
        mem[21] = 6'h3e;
        mem[22] = 6'h09;
        mem[23] = 6'h18;
        mem[24] = 6'h2e;
        mem[25] = 6'h01;
        mem[26] = 6'h33;
        mem[27] = 6'h11;
        mem[28] = 6'h07;
        mem[29] = 6'h3d;
        mem[30] = 6'h19;
        mem[31] = 6'h06;
        mem[32] = 6'h37;
        mem[33] = 6'h02;
        mem[34] = 6'h17;
        mem[35] = 6'h36;
        mem[36] = 6'h13;
        mem[37] = 6'h00;
        mem[38] = 6'h24;
        mem[39] = 6'h2b;
        mem[40] = 6'h2f;
        mem[41] = 6'h08;
        mem[42] = 6'h0e;
        mem[43] = 6'h0a;
        mem[44] = 6'h2c;
        mem[45] = 6'h15;
        mem[46] = 6'h31;
        mem[47] = 6'h27;
        mem[48] = 6'h1c;
        mem[49] = 6'h35;
        mem[50] = 6'h3a;
        mem[51] = 6'h26;
        mem[52] = 6'h32;
        mem[53] = 6'h23;
        mem[54] = 6'h2d;
        mem[55] = 6'h16;
        mem[56] = 6'h3f;
        mem[57] = 6'h12;
        mem[58] = 6'h0c;
        mem[59] = 6'h05;
        mem[60] = 6'h0b;
        mem[61] = 6'h20;
        mem[62] = 6'h21;
        mem[63] = 6'h1a;
    end
endmodule

module odo_sbox_small22(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h34;
        mem[1] = 6'h26;
        mem[2] = 6'h0c;
        mem[3] = 6'h1a;
        mem[4] = 6'h0e;
        mem[5] = 6'h1d;
        mem[6] = 6'h38;
        mem[7] = 6'h3d;
        mem[8] = 6'h35;
        mem[9] = 6'h21;
        mem[10] = 6'h1c;
        mem[11] = 6'h00;
        mem[12] = 6'h01;
        mem[13] = 6'h08;
        mem[14] = 6'h3b;
        mem[15] = 6'h1f;
        mem[16] = 6'h22;
        mem[17] = 6'h2c;
        mem[18] = 6'h15;
        mem[19] = 6'h2e;
        mem[20] = 6'h04;
        mem[21] = 6'h06;
        mem[22] = 6'h20;
        mem[23] = 6'h1e;
        mem[24] = 6'h10;
        mem[25] = 6'h09;
        mem[26] = 6'h37;
        mem[27] = 6'h31;
        mem[28] = 6'h14;
        mem[29] = 6'h0f;
        mem[30] = 6'h32;
        mem[31] = 6'h2a;
        mem[32] = 6'h33;
        mem[33] = 6'h24;
        mem[34] = 6'h3a;
        mem[35] = 6'h29;
        mem[36] = 6'h2f;
        mem[37] = 6'h3f;
        mem[38] = 6'h28;
        mem[39] = 6'h2b;
        mem[40] = 6'h02;
        mem[41] = 6'h1b;
        mem[42] = 6'h0d;
        mem[43] = 6'h25;
        mem[44] = 6'h23;
        mem[45] = 6'h19;
        mem[46] = 6'h0b;
        mem[47] = 6'h16;
        mem[48] = 6'h18;
        mem[49] = 6'h27;
        mem[50] = 6'h3c;
        mem[51] = 6'h36;
        mem[52] = 6'h03;
        mem[53] = 6'h39;
        mem[54] = 6'h30;
        mem[55] = 6'h07;
        mem[56] = 6'h17;
        mem[57] = 6'h05;
        mem[58] = 6'h12;
        mem[59] = 6'h11;
        mem[60] = 6'h3e;
        mem[61] = 6'h13;
        mem[62] = 6'h0a;
        mem[63] = 6'h2d;
    end
endmodule

module odo_sbox_small23(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h25;
        mem[1] = 6'h32;
        mem[2] = 6'h14;
        mem[3] = 6'h2e;
        mem[4] = 6'h29;
        mem[5] = 6'h0d;
        mem[6] = 6'h0a;
        mem[7] = 6'h15;
        mem[8] = 6'h26;
        mem[9] = 6'h0e;
        mem[10] = 6'h13;
        mem[11] = 6'h21;
        mem[12] = 6'h17;
        mem[13] = 6'h28;
        mem[14] = 6'h19;
        mem[15] = 6'h3b;
        mem[16] = 6'h23;
        mem[17] = 6'h39;
        mem[18] = 6'h22;
        mem[19] = 6'h38;
        mem[20] = 6'h2a;
        mem[21] = 6'h16;
        mem[22] = 6'h2b;
        mem[23] = 6'h3c;
        mem[24] = 6'h10;
        mem[25] = 6'h0f;
        mem[26] = 6'h31;
        mem[27] = 6'h3f;
        mem[28] = 6'h03;
        mem[29] = 6'h18;
        mem[30] = 6'h24;
        mem[31] = 6'h09;
        mem[32] = 6'h11;
        mem[33] = 6'h04;
        mem[34] = 6'h2f;
        mem[35] = 6'h1c;
        mem[36] = 6'h36;
        mem[37] = 6'h1f;
        mem[38] = 6'h3d;
        mem[39] = 6'h3e;
        mem[40] = 6'h33;
        mem[41] = 6'h35;
        mem[42] = 6'h30;
        mem[43] = 6'h02;
        mem[44] = 6'h3a;
        mem[45] = 6'h37;
        mem[46] = 6'h2d;
        mem[47] = 6'h1e;
        mem[48] = 6'h0c;
        mem[49] = 6'h2c;
        mem[50] = 6'h08;
        mem[51] = 6'h34;
        mem[52] = 6'h1b;
        mem[53] = 6'h06;
        mem[54] = 6'h07;
        mem[55] = 6'h12;
        mem[56] = 6'h05;
        mem[57] = 6'h20;
        mem[58] = 6'h00;
        mem[59] = 6'h01;
        mem[60] = 6'h27;
        mem[61] = 6'h1a;
        mem[62] = 6'h0b;
        mem[63] = 6'h1d;
    end
endmodule

module odo_sbox_small24(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0f;
        mem[1] = 6'h33;
        mem[2] = 6'h1a;
        mem[3] = 6'h27;
        mem[4] = 6'h20;
        mem[5] = 6'h19;
        mem[6] = 6'h09;
        mem[7] = 6'h1f;
        mem[8] = 6'h0c;
        mem[9] = 6'h02;
        mem[10] = 6'h39;
        mem[11] = 6'h3b;
        mem[12] = 6'h21;
        mem[13] = 6'h18;
        mem[14] = 6'h17;
        mem[15] = 6'h12;
        mem[16] = 6'h0b;
        mem[17] = 6'h2f;
        mem[18] = 6'h03;
        mem[19] = 6'h2d;
        mem[20] = 6'h1c;
        mem[21] = 6'h1e;
        mem[22] = 6'h04;
        mem[23] = 6'h2a;
        mem[24] = 6'h16;
        mem[25] = 6'h24;
        mem[26] = 6'h2b;
        mem[27] = 6'h15;
        mem[28] = 6'h00;
        mem[29] = 6'h1d;
        mem[30] = 6'h06;
        mem[31] = 6'h2c;
        mem[32] = 6'h07;
        mem[33] = 6'h3e;
        mem[34] = 6'h35;
        mem[35] = 6'h3f;
        mem[36] = 6'h36;
        mem[37] = 6'h25;
        mem[38] = 6'h11;
        mem[39] = 6'h05;
        mem[40] = 6'h1b;
        mem[41] = 6'h3c;
        mem[42] = 6'h3a;
        mem[43] = 6'h0e;
        mem[44] = 6'h30;
        mem[45] = 6'h28;
        mem[46] = 6'h13;
        mem[47] = 6'h34;
        mem[48] = 6'h08;
        mem[49] = 6'h26;
        mem[50] = 6'h10;
        mem[51] = 6'h22;
        mem[52] = 6'h29;
        mem[53] = 6'h37;
        mem[54] = 6'h23;
        mem[55] = 6'h01;
        mem[56] = 6'h31;
        mem[57] = 6'h2e;
        mem[58] = 6'h3d;
        mem[59] = 6'h0a;
        mem[60] = 6'h38;
        mem[61] = 6'h32;
        mem[62] = 6'h14;
        mem[63] = 6'h0d;
    end
endmodule

module odo_sbox_small25(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h36;
        mem[1] = 6'h14;
        mem[2] = 6'h19;
        mem[3] = 6'h2f;
        mem[4] = 6'h1a;
        mem[5] = 6'h1b;
        mem[6] = 6'h2b;
        mem[7] = 6'h0f;
        mem[8] = 6'h09;
        mem[9] = 6'h37;
        mem[10] = 6'h28;
        mem[11] = 6'h20;
        mem[12] = 6'h3e;
        mem[13] = 6'h27;
        mem[14] = 6'h04;
        mem[15] = 6'h29;
        mem[16] = 6'h35;
        mem[17] = 6'h22;
        mem[18] = 6'h21;
        mem[19] = 6'h06;
        mem[20] = 6'h0a;
        mem[21] = 6'h34;
        mem[22] = 6'h25;
        mem[23] = 6'h08;
        mem[24] = 6'h38;
        mem[25] = 6'h26;
        mem[26] = 6'h3b;
        mem[27] = 6'h3f;
        mem[28] = 6'h2d;
        mem[29] = 6'h3c;
        mem[30] = 6'h10;
        mem[31] = 6'h2a;
        mem[32] = 6'h15;
        mem[33] = 6'h1d;
        mem[34] = 6'h0d;
        mem[35] = 6'h11;
        mem[36] = 6'h33;
        mem[37] = 6'h30;
        mem[38] = 6'h07;
        mem[39] = 6'h0e;
        mem[40] = 6'h3d;
        mem[41] = 6'h2e;
        mem[42] = 6'h01;
        mem[43] = 6'h13;
        mem[44] = 6'h1e;
        mem[45] = 6'h24;
        mem[46] = 6'h23;
        mem[47] = 6'h31;
        mem[48] = 6'h39;
        mem[49] = 6'h02;
        mem[50] = 6'h16;
        mem[51] = 6'h18;
        mem[52] = 6'h12;
        mem[53] = 6'h2c;
        mem[54] = 6'h17;
        mem[55] = 6'h00;
        mem[56] = 6'h1f;
        mem[57] = 6'h3a;
        mem[58] = 6'h0b;
        mem[59] = 6'h05;
        mem[60] = 6'h1c;
        mem[61] = 6'h32;
        mem[62] = 6'h0c;
        mem[63] = 6'h03;
    end
endmodule

module odo_sbox_small26(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h08;
        mem[1] = 6'h03;
        mem[2] = 6'h39;
        mem[3] = 6'h38;
        mem[4] = 6'h20;
        mem[5] = 6'h30;
        mem[6] = 6'h31;
        mem[7] = 6'h24;
        mem[8] = 6'h25;
        mem[9] = 6'h06;
        mem[10] = 6'h05;
        mem[11] = 6'h2c;
        mem[12] = 6'h3a;
        mem[13] = 6'h16;
        mem[14] = 6'h13;
        mem[15] = 6'h1c;
        mem[16] = 6'h0d;
        mem[17] = 6'h34;
        mem[18] = 6'h01;
        mem[19] = 6'h3d;
        mem[20] = 6'h32;
        mem[21] = 6'h17;
        mem[22] = 6'h15;
        mem[23] = 6'h23;
        mem[24] = 6'h37;
        mem[25] = 6'h22;
        mem[26] = 6'h0c;
        mem[27] = 6'h26;
        mem[28] = 6'h28;
        mem[29] = 6'h3e;
        mem[30] = 6'h3c;
        mem[31] = 6'h2a;
        mem[32] = 6'h3b;
        mem[33] = 6'h21;
        mem[34] = 6'h1a;
        mem[35] = 6'h09;
        mem[36] = 6'h0b;
        mem[37] = 6'h35;
        mem[38] = 6'h2e;
        mem[39] = 6'h0e;
        mem[40] = 6'h18;
        mem[41] = 6'h10;
        mem[42] = 6'h27;
        mem[43] = 6'h0a;
        mem[44] = 6'h12;
        mem[45] = 6'h33;
        mem[46] = 6'h11;
        mem[47] = 6'h19;
        mem[48] = 6'h04;
        mem[49] = 6'h2f;
        mem[50] = 6'h29;
        mem[51] = 6'h1f;
        mem[52] = 6'h1e;
        mem[53] = 6'h1b;
        mem[54] = 6'h0f;
        mem[55] = 6'h2b;
        mem[56] = 6'h07;
        mem[57] = 6'h02;
        mem[58] = 6'h00;
        mem[59] = 6'h14;
        mem[60] = 6'h1d;
        mem[61] = 6'h36;
        mem[62] = 6'h3f;
        mem[63] = 6'h2d;
    end
endmodule

module odo_sbox_small27(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h12;
        mem[1] = 6'h02;
        mem[2] = 6'h09;
        mem[3] = 6'h3f;
        mem[4] = 6'h27;
        mem[5] = 6'h00;
        mem[6] = 6'h0c;
        mem[7] = 6'h2d;
        mem[8] = 6'h19;
        mem[9] = 6'h0b;
        mem[10] = 6'h37;
        mem[11] = 6'h2a;
        mem[12] = 6'h31;
        mem[13] = 6'h33;
        mem[14] = 6'h23;
        mem[15] = 6'h39;
        mem[16] = 6'h35;
        mem[17] = 6'h11;
        mem[18] = 6'h14;
        mem[19] = 6'h1e;
        mem[20] = 6'h03;
        mem[21] = 6'h1c;
        mem[22] = 6'h24;
        mem[23] = 6'h3c;
        mem[24] = 6'h3b;
        mem[25] = 6'h32;
        mem[26] = 6'h16;
        mem[27] = 6'h2f;
        mem[28] = 6'h0a;
        mem[29] = 6'h21;
        mem[30] = 6'h0f;
        mem[31] = 6'h1f;
        mem[32] = 6'h30;
        mem[33] = 6'h0d;
        mem[34] = 6'h04;
        mem[35] = 6'h2b;
        mem[36] = 6'h36;
        mem[37] = 6'h2c;
        mem[38] = 6'h06;
        mem[39] = 6'h13;
        mem[40] = 6'h38;
        mem[41] = 6'h15;
        mem[42] = 6'h3e;
        mem[43] = 6'h1d;
        mem[44] = 6'h2e;
        mem[45] = 6'h1a;
        mem[46] = 6'h10;
        mem[47] = 6'h3a;
        mem[48] = 6'h1b;
        mem[49] = 6'h22;
        mem[50] = 6'h17;
        mem[51] = 6'h25;
        mem[52] = 6'h34;
        mem[53] = 6'h20;
        mem[54] = 6'h0e;
        mem[55] = 6'h07;
        mem[56] = 6'h05;
        mem[57] = 6'h29;
        mem[58] = 6'h18;
        mem[59] = 6'h01;
        mem[60] = 6'h28;
        mem[61] = 6'h08;
        mem[62] = 6'h26;
        mem[63] = 6'h3d;
    end
endmodule

module odo_sbox_small28(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3a;
        mem[1] = 6'h17;
        mem[2] = 6'h0e;
        mem[3] = 6'h12;
        mem[4] = 6'h10;
        mem[5] = 6'h05;
        mem[6] = 6'h19;
        mem[7] = 6'h1d;
        mem[8] = 6'h14;
        mem[9] = 6'h0a;
        mem[10] = 6'h2a;
        mem[11] = 6'h38;
        mem[12] = 6'h0d;
        mem[13] = 6'h2b;
        mem[14] = 6'h34;
        mem[15] = 6'h0b;
        mem[16] = 6'h35;
        mem[17] = 6'h0c;
        mem[18] = 6'h18;
        mem[19] = 6'h1c;
        mem[20] = 6'h2e;
        mem[21] = 6'h0f;
        mem[22] = 6'h21;
        mem[23] = 6'h07;
        mem[24] = 6'h2f;
        mem[25] = 6'h27;
        mem[26] = 6'h00;
        mem[27] = 6'h24;
        mem[28] = 6'h20;
        mem[29] = 6'h26;
        mem[30] = 6'h04;
        mem[31] = 6'h31;
        mem[32] = 6'h02;
        mem[33] = 6'h1b;
        mem[34] = 6'h39;
        mem[35] = 6'h15;
        mem[36] = 6'h16;
        mem[37] = 6'h3d;
        mem[38] = 6'h09;
        mem[39] = 6'h01;
        mem[40] = 6'h29;
        mem[41] = 6'h3c;
        mem[42] = 6'h32;
        mem[43] = 6'h11;
        mem[44] = 6'h23;
        mem[45] = 6'h36;
        mem[46] = 6'h3b;
        mem[47] = 6'h06;
        mem[48] = 6'h13;
        mem[49] = 6'h03;
        mem[50] = 6'h25;
        mem[51] = 6'h33;
        mem[52] = 6'h1e;
        mem[53] = 6'h2c;
        mem[54] = 6'h08;
        mem[55] = 6'h37;
        mem[56] = 6'h1a;
        mem[57] = 6'h22;
        mem[58] = 6'h3f;
        mem[59] = 6'h1f;
        mem[60] = 6'h30;
        mem[61] = 6'h28;
        mem[62] = 6'h2d;
        mem[63] = 6'h3e;
    end
endmodule

module odo_sbox_small29(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1c;
        mem[1] = 6'h00;
        mem[2] = 6'h2e;
        mem[3] = 6'h23;
        mem[4] = 6'h08;
        mem[5] = 6'h18;
        mem[6] = 6'h3c;
        mem[7] = 6'h37;
        mem[8] = 6'h0e;
        mem[9] = 6'h06;
        mem[10] = 6'h3b;
        mem[11] = 6'h35;
        mem[12] = 6'h26;
        mem[13] = 6'h28;
        mem[14] = 6'h0a;
        mem[15] = 6'h09;
        mem[16] = 6'h1d;
        mem[17] = 6'h0d;
        mem[18] = 6'h17;
        mem[19] = 6'h36;
        mem[20] = 6'h2c;
        mem[21] = 6'h1e;
        mem[22] = 6'h2d;
        mem[23] = 6'h25;
        mem[24] = 6'h19;
        mem[25] = 6'h1b;
        mem[26] = 6'h2a;
        mem[27] = 6'h30;
        mem[28] = 6'h05;
        mem[29] = 6'h24;
        mem[30] = 6'h3f;
        mem[31] = 6'h14;
        mem[32] = 6'h34;
        mem[33] = 6'h33;
        mem[34] = 6'h32;
        mem[35] = 6'h12;
        mem[36] = 6'h10;
        mem[37] = 6'h31;
        mem[38] = 6'h0b;
        mem[39] = 6'h07;
        mem[40] = 6'h1f;
        mem[41] = 6'h21;
        mem[42] = 6'h13;
        mem[43] = 6'h20;
        mem[44] = 6'h0c;
        mem[45] = 6'h3e;
        mem[46] = 6'h2b;
        mem[47] = 6'h2f;
        mem[48] = 6'h15;
        mem[49] = 6'h1a;
        mem[50] = 6'h3d;
        mem[51] = 6'h0f;
        mem[52] = 6'h03;
        mem[53] = 6'h27;
        mem[54] = 6'h11;
        mem[55] = 6'h38;
        mem[56] = 6'h39;
        mem[57] = 6'h16;
        mem[58] = 6'h04;
        mem[59] = 6'h29;
        mem[60] = 6'h02;
        mem[61] = 6'h01;
        mem[62] = 6'h3a;
        mem[63] = 6'h22;
    end
endmodule

module odo_sbox_small30(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0a;
        mem[1] = 6'h06;
        mem[2] = 6'h1c;
        mem[3] = 6'h3b;
        mem[4] = 6'h34;
        mem[5] = 6'h10;
        mem[6] = 6'h30;
        mem[7] = 6'h15;
        mem[8] = 6'h2f;
        mem[9] = 6'h09;
        mem[10] = 6'h1a;
        mem[11] = 6'h25;
        mem[12] = 6'h22;
        mem[13] = 6'h14;
        mem[14] = 6'h27;
        mem[15] = 6'h31;
        mem[16] = 6'h33;
        mem[17] = 6'h3c;
        mem[18] = 6'h32;
        mem[19] = 6'h1d;
        mem[20] = 6'h17;
        mem[21] = 6'h36;
        mem[22] = 6'h3a;
        mem[23] = 6'h05;
        mem[24] = 6'h0c;
        mem[25] = 6'h0d;
        mem[26] = 6'h3d;
        mem[27] = 6'h3e;
        mem[28] = 6'h1f;
        mem[29] = 6'h12;
        mem[30] = 6'h28;
        mem[31] = 6'h23;
        mem[32] = 6'h26;
        mem[33] = 6'h11;
        mem[34] = 6'h2c;
        mem[35] = 6'h2d;
        mem[36] = 6'h0f;
        mem[37] = 6'h21;
        mem[38] = 6'h16;
        mem[39] = 6'h20;
        mem[40] = 6'h37;
        mem[41] = 6'h18;
        mem[42] = 6'h03;
        mem[43] = 6'h02;
        mem[44] = 6'h39;
        mem[45] = 6'h38;
        mem[46] = 6'h35;
        mem[47] = 6'h1b;
        mem[48] = 6'h2e;
        mem[49] = 6'h04;
        mem[50] = 6'h07;
        mem[51] = 6'h08;
        mem[52] = 6'h2a;
        mem[53] = 6'h00;
        mem[54] = 6'h0e;
        mem[55] = 6'h3f;
        mem[56] = 6'h01;
        mem[57] = 6'h29;
        mem[58] = 6'h19;
        mem[59] = 6'h1e;
        mem[60] = 6'h2b;
        mem[61] = 6'h0b;
        mem[62] = 6'h13;
        mem[63] = 6'h24;
    end
endmodule

module odo_sbox_small31(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h08;
        mem[1] = 6'h0b;
        mem[2] = 6'h1b;
        mem[3] = 6'h2c;
        mem[4] = 6'h32;
        mem[5] = 6'h00;
        mem[6] = 6'h15;
        mem[7] = 6'h24;
        mem[8] = 6'h2f;
        mem[9] = 6'h3d;
        mem[10] = 6'h14;
        mem[11] = 6'h38;
        mem[12] = 6'h1e;
        mem[13] = 6'h33;
        mem[14] = 6'h27;
        mem[15] = 6'h37;
        mem[16] = 6'h11;
        mem[17] = 6'h0f;
        mem[18] = 6'h0a;
        mem[19] = 6'h13;
        mem[20] = 6'h3f;
        mem[21] = 6'h1f;
        mem[22] = 6'h17;
        mem[23] = 6'h03;
        mem[24] = 6'h21;
        mem[25] = 6'h10;
        mem[26] = 6'h0e;
        mem[27] = 6'h3c;
        mem[28] = 6'h09;
        mem[29] = 6'h04;
        mem[30] = 6'h12;
        mem[31] = 6'h19;
        mem[32] = 6'h2d;
        mem[33] = 6'h39;
        mem[34] = 6'h02;
        mem[35] = 6'h1d;
        mem[36] = 6'h0c;
        mem[37] = 6'h29;
        mem[38] = 6'h28;
        mem[39] = 6'h3a;
        mem[40] = 6'h18;
        mem[41] = 6'h2a;
        mem[42] = 6'h26;
        mem[43] = 6'h23;
        mem[44] = 6'h2b;
        mem[45] = 6'h3b;
        mem[46] = 6'h1c;
        mem[47] = 6'h25;
        mem[48] = 6'h35;
        mem[49] = 6'h0d;
        mem[50] = 6'h30;
        mem[51] = 6'h1a;
        mem[52] = 6'h22;
        mem[53] = 6'h06;
        mem[54] = 6'h34;
        mem[55] = 6'h20;
        mem[56] = 6'h05;
        mem[57] = 6'h36;
        mem[58] = 6'h07;
        mem[59] = 6'h31;
        mem[60] = 6'h01;
        mem[61] = 6'h16;
        mem[62] = 6'h2e;
        mem[63] = 6'h3e;
    end
endmodule

module odo_sbox_small32(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0f;
        mem[1] = 6'h1a;
        mem[2] = 6'h02;
        mem[3] = 6'h21;
        mem[4] = 6'h1e;
        mem[5] = 6'h3f;
        mem[6] = 6'h2f;
        mem[7] = 6'h1c;
        mem[8] = 6'h26;
        mem[9] = 6'h0b;
        mem[10] = 6'h15;
        mem[11] = 6'h0e;
        mem[12] = 6'h25;
        mem[13] = 6'h14;
        mem[14] = 6'h19;
        mem[15] = 6'h23;
        mem[16] = 6'h0d;
        mem[17] = 6'h2d;
        mem[18] = 6'h36;
        mem[19] = 6'h1f;
        mem[20] = 6'h22;
        mem[21] = 6'h09;
        mem[22] = 6'h0c;
        mem[23] = 6'h24;
        mem[24] = 6'h04;
        mem[25] = 6'h32;
        mem[26] = 6'h29;
        mem[27] = 6'h17;
        mem[28] = 6'h35;
        mem[29] = 6'h2a;
        mem[30] = 6'h34;
        mem[31] = 6'h20;
        mem[32] = 6'h27;
        mem[33] = 6'h3c;
        mem[34] = 6'h2b;
        mem[35] = 6'h10;
        mem[36] = 6'h07;
        mem[37] = 6'h37;
        mem[38] = 6'h3d;
        mem[39] = 6'h00;
        mem[40] = 6'h2c;
        mem[41] = 6'h08;
        mem[42] = 6'h16;
        mem[43] = 6'h1d;
        mem[44] = 6'h31;
        mem[45] = 6'h39;
        mem[46] = 6'h30;
        mem[47] = 6'h2e;
        mem[48] = 6'h3e;
        mem[49] = 6'h03;
        mem[50] = 6'h0a;
        mem[51] = 6'h12;
        mem[52] = 6'h01;
        mem[53] = 6'h05;
        mem[54] = 6'h06;
        mem[55] = 6'h3b;
        mem[56] = 6'h13;
        mem[57] = 6'h3a;
        mem[58] = 6'h11;
        mem[59] = 6'h28;
        mem[60] = 6'h18;
        mem[61] = 6'h1b;
        mem[62] = 6'h33;
        mem[63] = 6'h38;
    end
endmodule

module odo_sbox_small33(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h38;
        mem[1] = 6'h1c;
        mem[2] = 6'h06;
        mem[3] = 6'h01;
        mem[4] = 6'h1d;
        mem[5] = 6'h39;
        mem[6] = 6'h3e;
        mem[7] = 6'h0e;
        mem[8] = 6'h1f;
        mem[9] = 6'h10;
        mem[10] = 6'h2b;
        mem[11] = 6'h30;
        mem[12] = 6'h15;
        mem[13] = 6'h33;
        mem[14] = 6'h2f;
        mem[15] = 6'h26;
        mem[16] = 6'h08;
        mem[17] = 6'h32;
        mem[18] = 6'h2c;
        mem[19] = 6'h09;
        mem[20] = 6'h07;
        mem[21] = 6'h1a;
        mem[22] = 6'h13;
        mem[23] = 6'h23;
        mem[24] = 6'h12;
        mem[25] = 6'h3c;
        mem[26] = 6'h29;
        mem[27] = 6'h34;
        mem[28] = 6'h19;
        mem[29] = 6'h21;
        mem[30] = 6'h0a;
        mem[31] = 6'h22;
        mem[32] = 6'h25;
        mem[33] = 6'h0c;
        mem[34] = 6'h0d;
        mem[35] = 6'h2d;
        mem[36] = 6'h17;
        mem[37] = 6'h36;
        mem[38] = 6'h18;
        mem[39] = 6'h3d;
        mem[40] = 6'h1b;
        mem[41] = 6'h20;
        mem[42] = 6'h28;
        mem[43] = 6'h1e;
        mem[44] = 6'h3a;
        mem[45] = 6'h02;
        mem[46] = 6'h31;
        mem[47] = 6'h0b;
        mem[48] = 6'h3b;
        mem[49] = 6'h24;
        mem[50] = 6'h00;
        mem[51] = 6'h3f;
        mem[52] = 6'h35;
        mem[53] = 6'h11;
        mem[54] = 6'h14;
        mem[55] = 6'h2a;
        mem[56] = 6'h2e;
        mem[57] = 6'h0f;
        mem[58] = 6'h04;
        mem[59] = 6'h27;
        mem[60] = 6'h05;
        mem[61] = 6'h37;
        mem[62] = 6'h16;
        mem[63] = 6'h03;
    end
endmodule

module odo_sbox_small34(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h32;
        mem[1] = 6'h04;
        mem[2] = 6'h23;
        mem[3] = 6'h21;
        mem[4] = 6'h3f;
        mem[5] = 6'h2a;
        mem[6] = 6'h1a;
        mem[7] = 6'h3b;
        mem[8] = 6'h3c;
        mem[9] = 6'h06;
        mem[10] = 6'h27;
        mem[11] = 6'h2d;
        mem[12] = 6'h0b;
        mem[13] = 6'h09;
        mem[14] = 6'h38;
        mem[15] = 6'h1c;
        mem[16] = 6'h39;
        mem[17] = 6'h1b;
        mem[18] = 6'h10;
        mem[19] = 6'h28;
        mem[20] = 6'h3e;
        mem[21] = 6'h1d;
        mem[22] = 6'h0c;
        mem[23] = 6'h01;
        mem[24] = 6'h20;
        mem[25] = 6'h25;
        mem[26] = 6'h29;
        mem[27] = 6'h36;
        mem[28] = 6'h17;
        mem[29] = 6'h0a;
        mem[30] = 6'h22;
        mem[31] = 6'h0e;
        mem[32] = 6'h07;
        mem[33] = 6'h3d;
        mem[34] = 6'h13;
        mem[35] = 6'h02;
        mem[36] = 6'h2e;
        mem[37] = 6'h26;
        mem[38] = 6'h18;
        mem[39] = 6'h37;
        mem[40] = 6'h2c;
        mem[41] = 6'h08;
        mem[42] = 6'h14;
        mem[43] = 6'h34;
        mem[44] = 6'h31;
        mem[45] = 6'h19;
        mem[46] = 6'h2f;
        mem[47] = 6'h03;
        mem[48] = 6'h2b;
        mem[49] = 6'h05;
        mem[50] = 6'h15;
        mem[51] = 6'h11;
        mem[52] = 6'h16;
        mem[53] = 6'h3a;
        mem[54] = 6'h1e;
        mem[55] = 6'h24;
        mem[56] = 6'h0f;
        mem[57] = 6'h12;
        mem[58] = 6'h00;
        mem[59] = 6'h33;
        mem[60] = 6'h35;
        mem[61] = 6'h1f;
        mem[62] = 6'h30;
        mem[63] = 6'h0d;
    end
endmodule

module odo_sbox_small35(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1a;
        mem[1] = 6'h37;
        mem[2] = 6'h2a;
        mem[3] = 6'h29;
        mem[4] = 6'h30;
        mem[5] = 6'h03;
        mem[6] = 6'h1d;
        mem[7] = 6'h16;
        mem[8] = 6'h0c;
        mem[9] = 6'h00;
        mem[10] = 6'h39;
        mem[11] = 6'h35;
        mem[12] = 6'h2b;
        mem[13] = 6'h04;
        mem[14] = 6'h15;
        mem[15] = 6'h1c;
        mem[16] = 6'h13;
        mem[17] = 6'h14;
        mem[18] = 6'h22;
        mem[19] = 6'h02;
        mem[20] = 6'h05;
        mem[21] = 6'h0e;
        mem[22] = 6'h3e;
        mem[23] = 6'h2d;
        mem[24] = 6'h0a;
        mem[25] = 6'h2c;
        mem[26] = 6'h32;
        mem[27] = 6'h09;
        mem[28] = 6'h2f;
        mem[29] = 6'h36;
        mem[30] = 6'h06;
        mem[31] = 6'h17;
        mem[32] = 6'h28;
        mem[33] = 6'h1b;
        mem[34] = 6'h24;
        mem[35] = 6'h19;
        mem[36] = 6'h0d;
        mem[37] = 6'h12;
        mem[38] = 6'h21;
        mem[39] = 6'h1f;
        mem[40] = 6'h0f;
        mem[41] = 6'h20;
        mem[42] = 6'h3f;
        mem[43] = 6'h2e;
        mem[44] = 6'h11;
        mem[45] = 6'h26;
        mem[46] = 6'h01;
        mem[47] = 6'h3d;
        mem[48] = 6'h10;
        mem[49] = 6'h07;
        mem[50] = 6'h1e;
        mem[51] = 6'h27;
        mem[52] = 6'h3b;
        mem[53] = 6'h25;
        mem[54] = 6'h18;
        mem[55] = 6'h31;
        mem[56] = 6'h08;
        mem[57] = 6'h34;
        mem[58] = 6'h38;
        mem[59] = 6'h3c;
        mem[60] = 6'h23;
        mem[61] = 6'h0b;
        mem[62] = 6'h33;
        mem[63] = 6'h3a;
    end
endmodule

module odo_sbox_small36(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2d;
        mem[1] = 6'h0b;
        mem[2] = 6'h2f;
        mem[3] = 6'h30;
        mem[4] = 6'h23;
        mem[5] = 6'h3c;
        mem[6] = 6'h08;
        mem[7] = 6'h2a;
        mem[8] = 6'h15;
        mem[9] = 6'h00;
        mem[10] = 6'h1a;
        mem[11] = 6'h0a;
        mem[12] = 6'h06;
        mem[13] = 6'h11;
        mem[14] = 6'h1f;
        mem[15] = 6'h29;
        mem[16] = 6'h37;
        mem[17] = 6'h12;
        mem[18] = 6'h3a;
        mem[19] = 6'h0c;
        mem[20] = 6'h13;
        mem[21] = 6'h3f;
        mem[22] = 6'h24;
        mem[23] = 6'h1b;
        mem[24] = 6'h0f;
        mem[25] = 6'h35;
        mem[26] = 6'h26;
        mem[27] = 6'h34;
        mem[28] = 6'h2b;
        mem[29] = 6'h19;
        mem[30] = 6'h1d;
        mem[31] = 6'h22;
        mem[32] = 6'h2e;
        mem[33] = 6'h18;
        mem[34] = 6'h09;
        mem[35] = 6'h32;
        mem[36] = 6'h20;
        mem[37] = 6'h02;
        mem[38] = 6'h28;
        mem[39] = 6'h0e;
        mem[40] = 6'h36;
        mem[41] = 6'h05;
        mem[42] = 6'h3d;
        mem[43] = 6'h16;
        mem[44] = 6'h2c;
        mem[45] = 6'h03;
        mem[46] = 6'h1c;
        mem[47] = 6'h07;
        mem[48] = 6'h27;
        mem[49] = 6'h1e;
        mem[50] = 6'h3e;
        mem[51] = 6'h10;
        mem[52] = 6'h17;
        mem[53] = 6'h25;
        mem[54] = 6'h31;
        mem[55] = 6'h33;
        mem[56] = 6'h01;
        mem[57] = 6'h21;
        mem[58] = 6'h04;
        mem[59] = 6'h0d;
        mem[60] = 6'h14;
        mem[61] = 6'h38;
        mem[62] = 6'h3b;
        mem[63] = 6'h39;
    end
endmodule

module odo_sbox_small37(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h18;
        mem[1] = 6'h36;
        mem[2] = 6'h20;
        mem[3] = 6'h10;
        mem[4] = 6'h3b;
        mem[5] = 6'h12;
        mem[6] = 6'h06;
        mem[7] = 6'h3f;
        mem[8] = 6'h22;
        mem[9] = 6'h24;
        mem[10] = 6'h28;
        mem[11] = 6'h00;
        mem[12] = 6'h37;
        mem[13] = 6'h3d;
        mem[14] = 6'h1f;
        mem[15] = 6'h2a;
        mem[16] = 6'h21;
        mem[17] = 6'h1a;
        mem[18] = 6'h0d;
        mem[19] = 6'h3c;
        mem[20] = 6'h2c;
        mem[21] = 6'h0f;
        mem[22] = 6'h0a;
        mem[23] = 6'h0c;
        mem[24] = 6'h01;
        mem[25] = 6'h33;
        mem[26] = 6'h19;
        mem[27] = 6'h09;
        mem[28] = 6'h31;
        mem[29] = 6'h2f;
        mem[30] = 6'h03;
        mem[31] = 6'h1c;
        mem[32] = 6'h38;
        mem[33] = 6'h13;
        mem[34] = 6'h16;
        mem[35] = 6'h17;
        mem[36] = 6'h04;
        mem[37] = 6'h27;
        mem[38] = 6'h02;
        mem[39] = 6'h05;
        mem[40] = 6'h32;
        mem[41] = 6'h14;
        mem[42] = 6'h1e;
        mem[43] = 6'h0e;
        mem[44] = 6'h1d;
        mem[45] = 6'h34;
        mem[46] = 6'h2b;
        mem[47] = 6'h23;
        mem[48] = 6'h1b;
        mem[49] = 6'h2d;
        mem[50] = 6'h11;
        mem[51] = 6'h30;
        mem[52] = 6'h26;
        mem[53] = 6'h08;
        mem[54] = 6'h35;
        mem[55] = 6'h25;
        mem[56] = 6'h0b;
        mem[57] = 6'h29;
        mem[58] = 6'h15;
        mem[59] = 6'h3e;
        mem[60] = 6'h07;
        mem[61] = 6'h3a;
        mem[62] = 6'h39;
        mem[63] = 6'h2e;
    end
endmodule

module odo_sbox_small38(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h23;
        mem[1] = 6'h18;
        mem[2] = 6'h1e;
        mem[3] = 6'h0f;
        mem[4] = 6'h1b;
        mem[5] = 6'h09;
        mem[6] = 6'h0c;
        mem[7] = 6'h06;
        mem[8] = 6'h2e;
        mem[9] = 6'h3e;
        mem[10] = 6'h03;
        mem[11] = 6'h08;
        mem[12] = 6'h34;
        mem[13] = 6'h0e;
        mem[14] = 6'h05;
        mem[15] = 6'h13;
        mem[16] = 6'h20;
        mem[17] = 6'h3f;
        mem[18] = 6'h3d;
        mem[19] = 6'h2a;
        mem[20] = 6'h21;
        mem[21] = 6'h3a;
        mem[22] = 6'h29;
        mem[23] = 6'h26;
        mem[24] = 6'h27;
        mem[25] = 6'h36;
        mem[26] = 6'h12;
        mem[27] = 6'h31;
        mem[28] = 6'h39;
        mem[29] = 6'h22;
        mem[30] = 6'h2d;
        mem[31] = 6'h1f;
        mem[32] = 6'h1c;
        mem[33] = 6'h17;
        mem[34] = 6'h01;
        mem[35] = 6'h0d;
        mem[36] = 6'h1a;
        mem[37] = 6'h25;
        mem[38] = 6'h3b;
        mem[39] = 6'h19;
        mem[40] = 6'h32;
        mem[41] = 6'h14;
        mem[42] = 6'h2c;
        mem[43] = 6'h11;
        mem[44] = 6'h33;
        mem[45] = 6'h1d;
        mem[46] = 6'h07;
        mem[47] = 6'h24;
        mem[48] = 6'h38;
        mem[49] = 6'h2b;
        mem[50] = 6'h28;
        mem[51] = 6'h2f;
        mem[52] = 6'h02;
        mem[53] = 6'h0a;
        mem[54] = 6'h35;
        mem[55] = 6'h37;
        mem[56] = 6'h16;
        mem[57] = 6'h10;
        mem[58] = 6'h04;
        mem[59] = 6'h15;
        mem[60] = 6'h0b;
        mem[61] = 6'h3c;
        mem[62] = 6'h30;
        mem[63] = 6'h00;
    end
endmodule

module odo_sbox_small39(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3f;
        mem[1] = 6'h36;
        mem[2] = 6'h1e;
        mem[3] = 6'h12;
        mem[4] = 6'h05;
        mem[5] = 6'h3a;
        mem[6] = 6'h2e;
        mem[7] = 6'h1c;
        mem[8] = 6'h25;
        mem[9] = 6'h35;
        mem[10] = 6'h3d;
        mem[11] = 6'h31;
        mem[12] = 6'h33;
        mem[13] = 6'h39;
        mem[14] = 6'h23;
        mem[15] = 6'h16;
        mem[16] = 6'h27;
        mem[17] = 6'h14;
        mem[18] = 6'h08;
        mem[19] = 6'h2a;
        mem[20] = 6'h38;
        mem[21] = 6'h1a;
        mem[22] = 6'h1f;
        mem[23] = 6'h2d;
        mem[24] = 6'h07;
        mem[25] = 6'h02;
        mem[26] = 6'h01;
        mem[27] = 6'h04;
        mem[28] = 6'h15;
        mem[29] = 6'h0c;
        mem[30] = 6'h2b;
        mem[31] = 6'h00;
        mem[32] = 6'h28;
        mem[33] = 6'h3c;
        mem[34] = 6'h1d;
        mem[35] = 6'h2f;
        mem[36] = 6'h2c;
        mem[37] = 6'h30;
        mem[38] = 6'h3b;
        mem[39] = 6'h1b;
        mem[40] = 6'h37;
        mem[41] = 6'h32;
        mem[42] = 6'h3e;
        mem[43] = 6'h22;
        mem[44] = 6'h29;
        mem[45] = 6'h24;
        mem[46] = 6'h09;
        mem[47] = 6'h18;
        mem[48] = 6'h10;
        mem[49] = 6'h19;
        mem[50] = 6'h20;
        mem[51] = 6'h13;
        mem[52] = 6'h03;
        mem[53] = 6'h26;
        mem[54] = 6'h0b;
        mem[55] = 6'h34;
        mem[56] = 6'h0d;
        mem[57] = 6'h0e;
        mem[58] = 6'h0a;
        mem[59] = 6'h0f;
        mem[60] = 6'h21;
        mem[61] = 6'h11;
        mem[62] = 6'h17;
        mem[63] = 6'h06;
    end
endmodule

module odo_sbox_large0(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    (* ram_style = "block" *) reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h2d0;
        mem[1] = 10'h35c;
        mem[2] = 10'h0e3;
        mem[3] = 10'h117;
        mem[4] = 10'h2fe;
        mem[5] = 10'h110;
        mem[6] = 10'h332;
        mem[7] = 10'h32d;
        mem[8] = 10'h380;
        mem[9] = 10'h382;
        mem[10] = 10'h018;
        mem[11] = 10'h374;
        mem[12] = 10'h23b;
        mem[13] = 10'h158;
        mem[14] = 10'h239;
        mem[15] = 10'h087;
        mem[16] = 10'h1a1;
        mem[17] = 10'h1d0;
        mem[18] = 10'h325;
        mem[19] = 10'h386;
        mem[20] = 10'h149;
        mem[21] = 10'h1a5;
        mem[22] = 10'h2bd;
        mem[23] = 10'h0ca;
        mem[24] = 10'h27a;
        mem[25] = 10'h2cc;
        mem[26] = 10'h031;
        mem[27] = 10'h135;
        mem[28] = 10'h2aa;
        mem[29] = 10'h2e1;
        mem[30] = 10'h24a;
        mem[31] = 10'h005;
        mem[32] = 10'h1c7;
        mem[33] = 10'h16e;
        mem[34] = 10'h3e7;
        mem[35] = 10'h0ed;
        mem[36] = 10'h137;
        mem[37] = 10'h0ad;
        mem[38] = 10'h320;
        mem[39] = 10'h28a;
        mem[40] = 10'h24c;
        mem[41] = 10'h283;
        mem[42] = 10'h0b0;
        mem[43] = 10'h048;
        mem[44] = 10'h0eb;
        mem[45] = 10'h153;
        mem[46] = 10'h217;
        mem[47] = 10'h12d;
        mem[48] = 10'h3c4;
        mem[49] = 10'h0cf;
        mem[50] = 10'h148;
        mem[51] = 10'h318;
        mem[52] = 10'h196;
        mem[53] = 10'h3f4;
        mem[54] = 10'h01b;
        mem[55] = 10'h3b5;
        mem[56] = 10'h04d;
        mem[57] = 10'h2f1;
        mem[58] = 10'h13c;
        mem[59] = 10'h28b;
        mem[60] = 10'h1c4;
        mem[61] = 10'h3c9;
        mem[62] = 10'h1f8;
        mem[63] = 10'h042;
        mem[64] = 10'h072;
        mem[65] = 10'h019;
        mem[66] = 10'h124;
        mem[67] = 10'h26e;
        mem[68] = 10'h09b;
        mem[69] = 10'h043;
        mem[70] = 10'h3b0;
        mem[71] = 10'h276;
        mem[72] = 10'h322;
        mem[73] = 10'h18f;
        mem[74] = 10'h0c3;
        mem[75] = 10'h308;
        mem[76] = 10'h17b;
        mem[77] = 10'h31d;
        mem[78] = 10'h3ba;
        mem[79] = 10'h28c;
        mem[80] = 10'h18e;
        mem[81] = 10'h3fa;
        mem[82] = 10'h2dc;
        mem[83] = 10'h0f9;
        mem[84] = 10'h314;
        mem[85] = 10'h21c;
        mem[86] = 10'h1ff;
        mem[87] = 10'h0e8;
        mem[88] = 10'h19d;
        mem[89] = 10'h3d3;
        mem[90] = 10'h22e;
        mem[91] = 10'h273;
        mem[92] = 10'h295;
        mem[93] = 10'h292;
        mem[94] = 10'h266;
        mem[95] = 10'h028;
        mem[96] = 10'h0cd;
        mem[97] = 10'h169;
        mem[98] = 10'h136;
        mem[99] = 10'h228;
        mem[100] = 10'h089;
        mem[101] = 10'h3d8;
        mem[102] = 10'h11a;
        mem[103] = 10'h253;
        mem[104] = 10'h1a9;
        mem[105] = 10'h0ee;
        mem[106] = 10'h077;
        mem[107] = 10'h209;
        mem[108] = 10'h0bc;
        mem[109] = 10'h2fa;
        mem[110] = 10'h398;
        mem[111] = 10'h2b7;
        mem[112] = 10'h24d;
        mem[113] = 10'h1f4;
        mem[114] = 10'h13a;
        mem[115] = 10'h342;
        mem[116] = 10'h202;
        mem[117] = 10'h24b;
        mem[118] = 10'h2b1;
        mem[119] = 10'h0ff;
        mem[120] = 10'h119;
        mem[121] = 10'h0db;
        mem[122] = 10'h3a0;
        mem[123] = 10'h0d7;
        mem[124] = 10'h0ab;
        mem[125] = 10'h192;
        mem[126] = 10'h354;
        mem[127] = 10'h161;
        mem[128] = 10'h2cf;
        mem[129] = 10'h10f;
        mem[130] = 10'h3b2;
        mem[131] = 10'h0d8;
        mem[132] = 10'h220;
        mem[133] = 10'h3e8;
        mem[134] = 10'h36e;
        mem[135] = 10'h376;
        mem[136] = 10'h306;
        mem[137] = 10'h3a8;
        mem[138] = 10'h358;
        mem[139] = 10'h01f;
        mem[140] = 10'h231;
        mem[141] = 10'h39f;
        mem[142] = 10'h33b;
        mem[143] = 10'h2de;
        mem[144] = 10'h19b;
        mem[145] = 10'h0aa;
        mem[146] = 10'h002;
        mem[147] = 10'h187;
        mem[148] = 10'h007;
        mem[149] = 10'h1e1;
        mem[150] = 10'h13e;
        mem[151] = 10'h13d;
        mem[152] = 10'h168;
        mem[153] = 10'h025;
        mem[154] = 10'h25a;
        mem[155] = 10'h2e3;
        mem[156] = 10'h2d7;
        mem[157] = 10'h267;
        mem[158] = 10'h38e;
        mem[159] = 10'h15b;
        mem[160] = 10'h21f;
        mem[161] = 10'h2ac;
        mem[162] = 10'h21d;
        mem[163] = 10'h256;
        mem[164] = 10'h262;
        mem[165] = 10'h05e;
        mem[166] = 10'h009;
        mem[167] = 10'h34e;
        mem[168] = 10'h26b;
        mem[169] = 10'h068;
        mem[170] = 10'h105;
        mem[171] = 10'h1e4;
        mem[172] = 10'h31e;
        mem[173] = 10'h112;
        mem[174] = 10'h272;
        mem[175] = 10'h170;
        mem[176] = 10'h194;
        mem[177] = 10'h235;
        mem[178] = 10'h200;
        mem[179] = 10'h33c;
        mem[180] = 10'h286;
        mem[181] = 10'h0fe;
        mem[182] = 10'h10d;
        mem[183] = 10'h3a7;
        mem[184] = 10'h02d;
        mem[185] = 10'h245;
        mem[186] = 10'h251;
        mem[187] = 10'h132;
        mem[188] = 10'h264;
        mem[189] = 10'h3f3;
        mem[190] = 10'h3be;
        mem[191] = 10'h1d6;
        mem[192] = 10'h27e;
        mem[193] = 10'h2ef;
        mem[194] = 10'h1b4;
        mem[195] = 10'h31f;
        mem[196] = 10'h39c;
        mem[197] = 10'h150;
        mem[198] = 10'h17d;
        mem[199] = 10'h02b;
        mem[200] = 10'h33a;
        mem[201] = 10'h1c3;
        mem[202] = 10'h115;
        mem[203] = 10'h2c3;
        mem[204] = 10'h249;
        mem[205] = 10'h017;
        mem[206] = 10'h257;
        mem[207] = 10'h229;
        mem[208] = 10'h2ce;
        mem[209] = 10'h29c;
        mem[210] = 10'h284;
        mem[211] = 10'h146;
        mem[212] = 10'h369;
        mem[213] = 10'h1cb;
        mem[214] = 10'h297;
        mem[215] = 10'h1b7;
        mem[216] = 10'h11f;
        mem[217] = 10'h1d7;
        mem[218] = 10'h1d1;
        mem[219] = 10'h28e;
        mem[220] = 10'h230;
        mem[221] = 10'h1c0;
        mem[222] = 10'h1fc;
        mem[223] = 10'h0c7;
        mem[224] = 10'h3aa;
        mem[225] = 10'h0e4;
        mem[226] = 10'h044;
        mem[227] = 10'h053;
        mem[228] = 10'h0bb;
        mem[229] = 10'h33f;
        mem[230] = 10'h299;
        mem[231] = 10'h316;
        mem[232] = 10'h34c;
        mem[233] = 10'h134;
        mem[234] = 10'h254;
        mem[235] = 10'h155;
        mem[236] = 10'h1ea;
        mem[237] = 10'h0fa;
        mem[238] = 10'h327;
        mem[239] = 10'h11e;
        mem[240] = 10'h1d8;
        mem[241] = 10'h23e;
        mem[242] = 10'h2e6;
        mem[243] = 10'h363;
        mem[244] = 10'h219;
        mem[245] = 10'h131;
        mem[246] = 10'h0bd;
        mem[247] = 10'h25b;
        mem[248] = 10'h07c;
        mem[249] = 10'h118;
        mem[250] = 10'h1ad;
        mem[251] = 10'h384;
        mem[252] = 10'h076;
        mem[253] = 10'h0e2;
        mem[254] = 10'h224;
        mem[255] = 10'h2e0;
        mem[256] = 10'h378;
        mem[257] = 10'h3db;
        mem[258] = 10'h31b;
        mem[259] = 10'h139;
        mem[260] = 10'h334;
        mem[261] = 10'h2ae;
        mem[262] = 10'h3b9;
        mem[263] = 10'h22f;
        mem[264] = 10'h1b3;
        mem[265] = 10'h213;
        mem[266] = 10'h0e6;
        mem[267] = 10'h2d5;
        mem[268] = 10'h2f2;
        mem[269] = 10'h091;
        mem[270] = 10'h3e0;
        mem[271] = 10'h387;
        mem[272] = 10'h22b;
        mem[273] = 10'h22d;
        mem[274] = 10'h1a2;
        mem[275] = 10'h107;
        mem[276] = 10'h03f;
        mem[277] = 10'h07a;
        mem[278] = 10'h191;
        mem[279] = 10'h3ca;
        mem[280] = 10'h157;
        mem[281] = 10'h29b;
        mem[282] = 10'h29e;
        mem[283] = 10'h06f;
        mem[284] = 10'h12b;
        mem[285] = 10'h309;
        mem[286] = 10'h06b;
        mem[287] = 10'h38b;
        mem[288] = 10'h159;
        mem[289] = 10'h3de;
        mem[290] = 10'h2eb;
        mem[291] = 10'h34f;
        mem[292] = 10'h09a;
        mem[293] = 10'h326;
        mem[294] = 10'h348;
        mem[295] = 10'h3c3;
        mem[296] = 10'h2a3;
        mem[297] = 10'h05c;
        mem[298] = 10'h3ef;
        mem[299] = 10'h294;
        mem[300] = 10'h179;
        mem[301] = 10'h057;
        mem[302] = 10'h35d;
        mem[303] = 10'h2af;
        mem[304] = 10'h2ba;
        mem[305] = 10'h0af;
        mem[306] = 10'h315;
        mem[307] = 10'h227;
        mem[308] = 10'h18b;
        mem[309] = 10'h0e9;
        mem[310] = 10'h289;
        mem[311] = 10'h081;
        mem[312] = 10'h2c0;
        mem[313] = 10'h23c;
        mem[314] = 10'h337;
        mem[315] = 10'h233;
        mem[316] = 10'h1ac;
        mem[317] = 10'h1a7;
        mem[318] = 10'h182;
        mem[319] = 10'h163;
        mem[320] = 10'h193;
        mem[321] = 10'h14d;
        mem[322] = 10'h2b4;
        mem[323] = 10'h30e;
        mem[324] = 10'h2da;
        mem[325] = 10'h27c;
        mem[326] = 10'h186;
        mem[327] = 10'h0c5;
        mem[328] = 10'h3df;
        mem[329] = 10'h3fc;
        mem[330] = 10'h3e5;
        mem[331] = 10'h1e7;
        mem[332] = 10'h238;
        mem[333] = 10'h0c1;
        mem[334] = 10'h28f;
        mem[335] = 10'h1df;
        mem[336] = 10'h1b1;
        mem[337] = 10'h102;
        mem[338] = 10'h2a9;
        mem[339] = 10'h21a;
        mem[340] = 10'h2d9;
        mem[341] = 10'h0fc;
        mem[342] = 10'h215;
        mem[343] = 10'h0a5;
        mem[344] = 10'h3ec;
        mem[345] = 10'h1d5;
        mem[346] = 10'h2f8;
        mem[347] = 10'h1b8;
        mem[348] = 10'h389;
        mem[349] = 10'h00d;
        mem[350] = 10'h25f;
        mem[351] = 10'h0e7;
        mem[352] = 10'h379;
        mem[353] = 10'h3a3;
        mem[354] = 10'h172;
        mem[355] = 10'h114;
        mem[356] = 10'h1fd;
        mem[357] = 10'h16c;
        mem[358] = 10'h29d;
        mem[359] = 10'h0b8;
        mem[360] = 10'h0ba;
        mem[361] = 10'h1c1;
        mem[362] = 10'h211;
        mem[363] = 10'h18d;
        mem[364] = 10'h3e4;
        mem[365] = 10'h0f3;
        mem[366] = 10'h244;
        mem[367] = 10'h023;
        mem[368] = 10'h321;
        mem[369] = 10'h0b5;
        mem[370] = 10'h10b;
        mem[371] = 10'h37b;
        mem[372] = 10'h36b;
        mem[373] = 10'h177;
        mem[374] = 10'h097;
        mem[375] = 10'h18a;
        mem[376] = 10'h255;
        mem[377] = 10'h083;
        mem[378] = 10'h261;
        mem[379] = 10'h22c;
        mem[380] = 10'h368;
        mem[381] = 10'h095;
        mem[382] = 10'h3f9;
        mem[383] = 10'h199;
        mem[384] = 10'h3c7;
        mem[385] = 10'h0a3;
        mem[386] = 10'h2a5;
        mem[387] = 10'h207;
        mem[388] = 10'h3b4;
        mem[389] = 10'h121;
        mem[390] = 10'h0b4;
        mem[391] = 10'h30c;
        mem[392] = 10'h00e;
        mem[393] = 10'h16d;
        mem[394] = 10'h180;
        mem[395] = 10'h37d;
        mem[396] = 10'h07f;
        mem[397] = 10'h1ec;
        mem[398] = 10'h34b;
        mem[399] = 10'h11c;
        mem[400] = 10'h130;
        mem[401] = 10'h301;
        mem[402] = 10'h069;
        mem[403] = 10'h285;
        mem[404] = 10'h205;
        mem[405] = 10'h252;
        mem[406] = 10'h2ee;
        mem[407] = 10'h3cc;
        mem[408] = 10'h1cd;
        mem[409] = 10'h373;
        mem[410] = 10'h399;
        mem[411] = 10'h12a;
        mem[412] = 10'h147;
        mem[413] = 10'h01c;
        mem[414] = 10'h0d6;
        mem[415] = 10'h3f6;
        mem[416] = 10'h0a8;
        mem[417] = 10'h080;
        mem[418] = 10'h39a;
        mem[419] = 10'h390;
        mem[420] = 10'h3ce;
        mem[421] = 10'h28d;
        mem[422] = 10'h2e9;
        mem[423] = 10'h324;
        mem[424] = 10'h10c;
        mem[425] = 10'h2b2;
        mem[426] = 10'h17f;
        mem[427] = 10'h000;
        mem[428] = 10'h19c;
        mem[429] = 10'h15f;
        mem[430] = 10'h01a;
        mem[431] = 10'h367;
        mem[432] = 10'h3d1;
        mem[433] = 10'h1e0;
        mem[434] = 10'h345;
        mem[435] = 10'h2f0;
        mem[436] = 10'h13f;
        mem[437] = 10'h11d;
        mem[438] = 10'h323;
        mem[439] = 10'h287;
        mem[440] = 10'h293;
        mem[441] = 10'h371;
        mem[442] = 10'h15d;
        mem[443] = 10'h17c;
        mem[444] = 10'h09d;
        mem[445] = 10'h24e;
        mem[446] = 10'h15c;
        mem[447] = 10'h060;
        mem[448] = 10'h246;
        mem[449] = 10'h30a;
        mem[450] = 10'h32b;
        mem[451] = 10'h0c4;
        mem[452] = 10'h2d4;
        mem[453] = 10'h3ac;
        mem[454] = 10'h2c5;
        mem[455] = 10'h26d;
        mem[456] = 10'h2fd;
        mem[457] = 10'h0ac;
        mem[458] = 10'h0cb;
        mem[459] = 10'h14e;
        mem[460] = 10'h078;
        mem[461] = 10'h0a6;
        mem[462] = 10'h0fd;
        mem[463] = 10'h14c;
        mem[464] = 10'h3cf;
        mem[465] = 10'h25c;
        mem[466] = 10'h26a;
        mem[467] = 10'h35e;
        mem[468] = 10'h02a;
        mem[469] = 10'h30d;
        mem[470] = 10'h0ef;
        mem[471] = 10'h0d2;
        mem[472] = 10'h388;
        mem[473] = 10'h39d;
        mem[474] = 10'h1e5;
        mem[475] = 10'h392;
        mem[476] = 10'h344;
        mem[477] = 10'h311;
        mem[478] = 10'h0c2;
        mem[479] = 10'h0a4;
        mem[480] = 10'h020;
        mem[481] = 10'h1b6;
        mem[482] = 10'h2db;
        mem[483] = 10'h222;
        mem[484] = 10'h218;
        mem[485] = 10'h2e5;
        mem[486] = 10'h2b5;
        mem[487] = 10'h383;
        mem[488] = 10'h012;
        mem[489] = 10'h288;
        mem[490] = 10'h1a6;
        mem[491] = 10'h17e;
        mem[492] = 10'h052;
        mem[493] = 10'h290;
        mem[494] = 10'h265;
        mem[495] = 10'h14b;
        mem[496] = 10'h2f9;
        mem[497] = 10'h1fa;
        mem[498] = 10'h055;
        mem[499] = 10'h041;
        mem[500] = 10'h2e8;
        mem[501] = 10'h3a5;
        mem[502] = 10'h385;
        mem[503] = 10'h3d7;
        mem[504] = 10'h021;
        mem[505] = 10'h2ed;
        mem[506] = 10'h352;
        mem[507] = 10'h2bb;
        mem[508] = 10'h0b6;
        mem[509] = 10'h04f;
        mem[510] = 10'h223;
        mem[511] = 10'h154;
        mem[512] = 10'h3f5;
        mem[513] = 10'h333;
        mem[514] = 10'h11b;
        mem[515] = 10'h3ae;
        mem[516] = 10'h397;
        mem[517] = 10'h2a4;
        mem[518] = 10'h079;
        mem[519] = 10'h1e6;
        mem[520] = 10'h0c9;
        mem[521] = 10'h258;
        mem[522] = 10'h07d;
        mem[523] = 10'h274;
        mem[524] = 10'h176;
        mem[525] = 10'h35b;
        mem[526] = 10'h16f;
        mem[527] = 10'h32e;
        mem[528] = 10'h206;
        mem[529] = 10'h22a;
        mem[530] = 10'h395;
        mem[531] = 10'h3b8;
        mem[532] = 10'h338;
        mem[533] = 10'h1ba;
        mem[534] = 10'h016;
        mem[535] = 10'h00c;
        mem[536] = 10'h1e3;
        mem[537] = 10'h008;
        mem[538] = 10'h305;
        mem[539] = 10'h116;
        mem[540] = 10'h280;
        mem[541] = 10'h103;
        mem[542] = 10'h3c0;
        mem[543] = 10'h34a;
        mem[544] = 10'h06c;
        mem[545] = 10'h123;
        mem[546] = 10'h1d2;
        mem[547] = 10'h33d;
        mem[548] = 10'h0d0;
        mem[549] = 10'h36a;
        mem[550] = 10'h355;
        mem[551] = 10'h040;
        mem[552] = 10'h3a9;
        mem[553] = 10'h36c;
        mem[554] = 10'h2c4;
        mem[555] = 10'h16b;
        mem[556] = 10'h2f5;
        mem[557] = 10'h2b3;
        mem[558] = 10'h152;
        mem[559] = 10'h188;
        mem[560] = 10'h34d;
        mem[561] = 10'h1ae;
        mem[562] = 10'h15e;
        mem[563] = 10'h058;
        mem[564] = 10'h3ea;
        mem[565] = 10'h08b;
        mem[566] = 10'h059;
        mem[567] = 10'h175;
        mem[568] = 10'h065;
        mem[569] = 10'h0f7;
        mem[570] = 10'h2b9;
        mem[571] = 10'h221;
        mem[572] = 10'h3c1;
        mem[573] = 10'h0f8;
        mem[574] = 10'h381;
        mem[575] = 10'h06d;
        mem[576] = 10'h3e6;
        mem[577] = 10'h1ca;
        mem[578] = 10'h09c;
        mem[579] = 10'h013;
        mem[580] = 10'h1e9;
        mem[581] = 10'h1ce;
        mem[582] = 10'h375;
        mem[583] = 10'h061;
        mem[584] = 10'h2d2;
        mem[585] = 10'h1f7;
        mem[586] = 10'h38a;
        mem[587] = 10'h08c;
        mem[588] = 10'h1bd;
        mem[589] = 10'h08a;
        mem[590] = 10'h15a;
        mem[591] = 10'h298;
        mem[592] = 10'h029;
        mem[593] = 10'h1bb;
        mem[594] = 10'h084;
        mem[595] = 10'h2e2;
        mem[596] = 10'h14a;
        mem[597] = 10'h09f;
        mem[598] = 10'h2c6;
        mem[599] = 10'h0b3;
        mem[600] = 10'h0ea;
        mem[601] = 10'h2ec;
        mem[602] = 10'h39b;
        mem[603] = 10'h35f;
        mem[604] = 10'h2c7;
        mem[605] = 10'h2c9;
        mem[606] = 10'h13b;
        mem[607] = 10'h198;
        mem[608] = 10'h304;
        mem[609] = 10'h03a;
        mem[610] = 10'h201;
        mem[611] = 10'h370;
        mem[612] = 10'h045;
        mem[613] = 10'h046;
        mem[614] = 10'h329;
        mem[615] = 10'h056;
        mem[616] = 10'h156;
        mem[617] = 10'h3cd;
        mem[618] = 10'h3ad;
        mem[619] = 10'h39e;
        mem[620] = 10'h0a2;
        mem[621] = 10'h195;
        mem[622] = 10'h2df;
        mem[623] = 10'h3f8;
        mem[624] = 10'h06a;
        mem[625] = 10'h1a0;
        mem[626] = 10'h086;
        mem[627] = 10'h071;
        mem[628] = 10'h3a2;
        mem[629] = 10'h162;
        mem[630] = 10'h04c;
        mem[631] = 10'h3e2;
        mem[632] = 10'h2b0;
        mem[633] = 10'h126;
        mem[634] = 10'h335;
        mem[635] = 10'h0df;
        mem[636] = 10'h3ee;
        mem[637] = 10'h259;
        mem[638] = 10'h0e1;
        mem[639] = 10'h075;
        mem[640] = 10'h1a4;
        mem[641] = 10'h02f;
        mem[642] = 10'h26c;
        mem[643] = 10'h038;
        mem[644] = 10'h00f;
        mem[645] = 10'h1ed;
        mem[646] = 10'h033;
        mem[647] = 10'h1c2;
        mem[648] = 10'h27d;
        mem[649] = 10'h23d;
        mem[650] = 10'h0c8;
        mem[651] = 10'h0e0;
        mem[652] = 10'h21b;
        mem[653] = 10'h06e;
        mem[654] = 10'h0f5;
        mem[655] = 10'h23a;
        mem[656] = 10'h3ff;
        mem[657] = 10'h03c;
        mem[658] = 10'h047;
        mem[659] = 10'h29a;
        mem[660] = 10'h275;
        mem[661] = 10'h1b9;
        mem[662] = 10'h066;
        mem[663] = 10'h20a;
        mem[664] = 10'h240;
        mem[665] = 10'h173;
        mem[666] = 10'h085;
        mem[667] = 10'h01e;
        mem[668] = 10'h2ca;
        mem[669] = 10'h279;
        mem[670] = 10'h0dc;
        mem[671] = 10'h015;
        mem[672] = 10'h330;
        mem[673] = 10'h1f1;
        mem[674] = 10'h241;
        mem[675] = 10'h1f9;
        mem[676] = 10'h0ae;
        mem[677] = 10'h032;
        mem[678] = 10'h0b1;
        mem[679] = 10'h3c8;
        mem[680] = 10'h3d4;
        mem[681] = 10'h291;
        mem[682] = 10'h022;
        mem[683] = 10'h32a;
        mem[684] = 10'h027;
        mem[685] = 10'h04b;
        mem[686] = 10'h099;
        mem[687] = 10'h2d3;
        mem[688] = 10'h011;
        mem[689] = 10'h341;
        mem[690] = 10'h3f7;
        mem[691] = 10'h31a;
        mem[692] = 10'h2bc;
        mem[693] = 10'h104;
        mem[694] = 10'h128;
        mem[695] = 10'h164;
        mem[696] = 10'h2a6;
        mem[697] = 10'h05d;
        mem[698] = 10'h1f2;
        mem[699] = 10'h208;
        mem[700] = 10'h003;
        mem[701] = 10'h339;
        mem[702] = 10'h037;
        mem[703] = 10'h20c;
        mem[704] = 10'h036;
        mem[705] = 10'h10e;
        mem[706] = 10'h05f;
        mem[707] = 10'h1dd;
        mem[708] = 10'h1ee;
        mem[709] = 10'h2d6;
        mem[710] = 10'h26f;
        mem[711] = 10'h141;
        mem[712] = 10'h250;
        mem[713] = 10'h226;
        mem[714] = 10'h1fe;
        mem[715] = 10'h1de;
        mem[716] = 10'h109;
        mem[717] = 10'h3ab;
        mem[718] = 10'h05b;
        mem[719] = 10'h20e;
        mem[720] = 10'h151;
        mem[721] = 10'h3cb;
        mem[722] = 10'h1c6;
        mem[723] = 10'h160;
        mem[724] = 10'h350;
        mem[725] = 10'h174;
        mem[726] = 10'h1f5;
        mem[727] = 10'h08f;
        mem[728] = 10'h1bf;
        mem[729] = 10'h396;
        mem[730] = 10'h185;
        mem[731] = 10'h101;
        mem[732] = 10'h100;
        mem[733] = 10'h351;
        mem[734] = 10'h2b6;
        mem[735] = 10'h03e;
        mem[736] = 10'h1b2;
        mem[737] = 10'h346;
        mem[738] = 10'h05a;
        mem[739] = 10'h319;
        mem[740] = 10'h24f;
        mem[741] = 10'h2cd;
        mem[742] = 10'h1aa;
        mem[743] = 10'h23f;
        mem[744] = 10'h122;
        mem[745] = 10'h296;
        mem[746] = 10'h0a9;
        mem[747] = 10'h178;
        mem[748] = 10'h2e4;
        mem[749] = 10'h3da;
        mem[750] = 10'h1e2;
        mem[751] = 10'h364;
        mem[752] = 10'h2ad;
        mem[753] = 10'h004;
        mem[754] = 10'h2fc;
        mem[755] = 10'h1b5;
        mem[756] = 10'h04a;
        mem[757] = 10'h353;
        mem[758] = 10'h145;
        mem[759] = 10'h210;
        mem[760] = 10'h2a7;
        mem[761] = 10'h19a;
        mem[762] = 10'h14f;
        mem[763] = 10'h2ff;
        mem[764] = 10'h225;
        mem[765] = 10'h38f;
        mem[766] = 10'h37c;
        mem[767] = 10'h31c;
        mem[768] = 10'h171;
        mem[769] = 10'h236;
        mem[770] = 10'h3d2;
        mem[771] = 10'h30b;
        mem[772] = 10'h3bf;
        mem[773] = 10'h377;
        mem[774] = 10'h1db;
        mem[775] = 10'h312;
        mem[776] = 10'h08e;
        mem[777] = 10'h391;
        mem[778] = 10'h0c0;
        mem[779] = 10'h0f4;
        mem[780] = 10'h357;
        mem[781] = 10'h073;
        mem[782] = 10'h096;
        mem[783] = 10'h1f6;
        mem[784] = 10'h1f3;
        mem[785] = 10'h064;
        mem[786] = 10'h12e;
        mem[787] = 10'h36f;
        mem[788] = 10'h3c2;
        mem[789] = 10'h232;
        mem[790] = 10'h37a;
        mem[791] = 10'h183;
        mem[792] = 10'h03b;
        mem[793] = 10'h074;
        mem[794] = 10'h0b2;
        mem[795] = 10'h366;
        mem[796] = 10'h38d;
        mem[797] = 10'h0fb;
        mem[798] = 10'h1d4;
        mem[799] = 10'h1e8;
        mem[800] = 10'h0d4;
        mem[801] = 10'h30f;
        mem[802] = 10'h3e1;
        mem[803] = 10'h1ab;
        mem[804] = 10'h02c;
        mem[805] = 10'h039;
        mem[806] = 10'h27f;
        mem[807] = 10'h2fb;
        mem[808] = 10'h035;
        mem[809] = 10'h0d5;
        mem[810] = 10'h0de;
        mem[811] = 10'h2bf;
        mem[812] = 10'h281;
        mem[813] = 10'h0a0;
        mem[814] = 10'h0ce;
        mem[815] = 10'h070;
        mem[816] = 10'h328;
        mem[817] = 10'h0c6;
        mem[818] = 10'h282;
        mem[819] = 10'h3b6;
        mem[820] = 10'h165;
        mem[821] = 10'h1b0;
        mem[822] = 10'h263;
        mem[823] = 10'h1a3;
        mem[824] = 10'h277;
        mem[825] = 10'h062;
        mem[826] = 10'h3f1;
        mem[827] = 10'h010;
        mem[828] = 10'h3d0;
        mem[829] = 10'h3e9;
        mem[830] = 10'h1cf;
        mem[831] = 10'h216;
        mem[832] = 10'h144;
        mem[833] = 10'h260;
        mem[834] = 10'h063;
        mem[835] = 10'h1da;
        mem[836] = 10'h3d5;
        mem[837] = 10'h268;
        mem[838] = 10'h1bc;
        mem[839] = 10'h204;
        mem[840] = 10'h35a;
        mem[841] = 10'h3bb;
        mem[842] = 10'h3a1;
        mem[843] = 10'h050;
        mem[844] = 10'h18c;
        mem[845] = 10'h133;
        mem[846] = 10'h1a8;
        mem[847] = 10'h108;
        mem[848] = 10'h0b9;
        mem[849] = 10'h1c5;
        mem[850] = 10'h37e;
        mem[851] = 10'h362;
        mem[852] = 10'h1c9;
        mem[853] = 10'h0d1;
        mem[854] = 10'h1cc;
        mem[855] = 10'h02e;
        mem[856] = 10'h140;
        mem[857] = 10'h0e5;
        mem[858] = 10'h166;
        mem[859] = 10'h313;
        mem[860] = 10'h09e;
        mem[861] = 10'h19f;
        mem[862] = 10'h03d;
        mem[863] = 10'h1fb;
        mem[864] = 10'h3e3;
        mem[865] = 10'h2b8;
        mem[866] = 10'h33e;
        mem[867] = 10'h051;
        mem[868] = 10'h1ef;
        mem[869] = 10'h127;
        mem[870] = 10'h0f0;
        mem[871] = 10'h2a0;
        mem[872] = 10'h3bd;
        mem[873] = 10'h093;
        mem[874] = 10'h2ab;
        mem[875] = 10'h120;
        mem[876] = 10'h2f4;
        mem[877] = 10'h19e;
        mem[878] = 10'h030;
        mem[879] = 10'h0da;
        mem[880] = 10'h106;
        mem[881] = 10'h248;
        mem[882] = 10'h0be;
        mem[883] = 10'h006;
        mem[884] = 10'h2d8;
        mem[885] = 10'h317;
        mem[886] = 10'h361;
        mem[887] = 10'h142;
        mem[888] = 10'h271;
        mem[889] = 10'h014;
        mem[890] = 10'h32c;
        mem[891] = 10'h349;
        mem[892] = 10'h0b7;
        mem[893] = 10'h0a1;
        mem[894] = 10'h049;
        mem[895] = 10'h27b;
        mem[896] = 10'h0dd;
        mem[897] = 10'h08d;
        mem[898] = 10'h3d9;
        mem[899] = 10'h3fb;
        mem[900] = 10'h2f7;
        mem[901] = 10'h3bc;
        mem[902] = 10'h1dc;
        mem[903] = 10'h37f;
        mem[904] = 10'h365;
        mem[905] = 10'h214;
        mem[906] = 10'h1be;
        mem[907] = 10'h2d1;
        mem[908] = 10'h2c2;
        mem[909] = 10'h302;
        mem[910] = 10'h343;
        mem[911] = 10'h190;
        mem[912] = 10'h234;
        mem[913] = 10'h310;
        mem[914] = 10'h1d9;
        mem[915] = 10'h300;
        mem[916] = 10'h197;
        mem[917] = 10'h2cb;
        mem[918] = 10'h2e7;
        mem[919] = 10'h2f3;
        mem[920] = 10'h2dd;
        mem[921] = 10'h0ec;
        mem[922] = 10'h094;
        mem[923] = 10'h1af;
        mem[924] = 10'h167;
        mem[925] = 10'h184;
        mem[926] = 10'h2a8;
        mem[927] = 10'h0f6;
        mem[928] = 10'h347;
        mem[929] = 10'h067;
        mem[930] = 10'h2be;
        mem[931] = 10'h247;
        mem[932] = 10'h242;
        mem[933] = 10'h36d;
        mem[934] = 10'h359;
        mem[935] = 10'h3b3;
        mem[936] = 10'h21e;
        mem[937] = 10'h269;
        mem[938] = 10'h10a;
        mem[939] = 10'h243;
        mem[940] = 10'h394;
        mem[941] = 10'h0d9;
        mem[942] = 10'h17a;
        mem[943] = 10'h0d3;
        mem[944] = 10'h3f0;
        mem[945] = 10'h3fd;
        mem[946] = 10'h356;
        mem[947] = 10'h2f6;
        mem[948] = 10'h3dd;
        mem[949] = 10'h125;
        mem[950] = 10'h237;
        mem[951] = 10'h393;
        mem[952] = 10'h1f0;
        mem[953] = 10'h3a6;
        mem[954] = 10'h3b1;
        mem[955] = 10'h203;
        mem[956] = 10'h32f;
        mem[957] = 10'h098;
        mem[958] = 10'h3a4;
        mem[959] = 10'h3dc;
        mem[960] = 10'h07e;
        mem[961] = 10'h336;
        mem[962] = 10'h138;
        mem[963] = 10'h034;
        mem[964] = 10'h307;
        mem[965] = 10'h12c;
        mem[966] = 10'h113;
        mem[967] = 10'h3f2;
        mem[968] = 10'h3b7;
        mem[969] = 10'h07b;
        mem[970] = 10'h2a2;
        mem[971] = 10'h270;
        mem[972] = 10'h340;
        mem[973] = 10'h2a1;
        mem[974] = 10'h088;
        mem[975] = 10'h20d;
        mem[976] = 10'h1eb;
        mem[977] = 10'h04e;
        mem[978] = 10'h01d;
        mem[979] = 10'h143;
        mem[980] = 10'h2ea;
        mem[981] = 10'h00a;
        mem[982] = 10'h3ed;
        mem[983] = 10'h3fe;
        mem[984] = 10'h054;
        mem[985] = 10'h360;
        mem[986] = 10'h372;
        mem[987] = 10'h0a7;
        mem[988] = 10'h189;
        mem[989] = 10'h25e;
        mem[990] = 10'h1c8;
        mem[991] = 10'h0cc;
        mem[992] = 10'h38c;
        mem[993] = 10'h3c6;
        mem[994] = 10'h0f2;
        mem[995] = 10'h2c8;
        mem[996] = 10'h111;
        mem[997] = 10'h090;
        mem[998] = 10'h16a;
        mem[999] = 10'h1d3;
        mem[1000] = 10'h092;
        mem[1001] = 10'h3d6;
        mem[1002] = 10'h212;
        mem[1003] = 10'h0f1;
        mem[1004] = 10'h3c5;
        mem[1005] = 10'h278;
        mem[1006] = 10'h0bf;
        mem[1007] = 10'h129;
        mem[1008] = 10'h181;
        mem[1009] = 10'h3af;
        mem[1010] = 10'h12f;
        mem[1011] = 10'h082;
        mem[1012] = 10'h001;
        mem[1013] = 10'h29f;
        mem[1014] = 10'h026;
        mem[1015] = 10'h3eb;
        mem[1016] = 10'h331;
        mem[1017] = 10'h00b;
        mem[1018] = 10'h25d;
        mem[1019] = 10'h20b;
        mem[1020] = 10'h024;
        mem[1021] = 10'h303;
        mem[1022] = 10'h20f;
        mem[1023] = 10'h2c1;
    end
endmodule

module odo_sbox_large1(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    (* ram_style = "block" *) reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h1dc;
        mem[1] = 10'h21e;
        mem[2] = 10'h325;
        mem[3] = 10'h329;
        mem[4] = 10'h042;
        mem[5] = 10'h16e;
        mem[6] = 10'h0dc;
        mem[7] = 10'h306;
        mem[8] = 10'h372;
        mem[9] = 10'h1e6;
        mem[10] = 10'h34e;
        mem[11] = 10'h1ea;
        mem[12] = 10'h132;
        mem[13] = 10'h379;
        mem[14] = 10'h07b;
        mem[15] = 10'h3a8;
        mem[16] = 10'h07f;
        mem[17] = 10'h1c9;
        mem[18] = 10'h00a;
        mem[19] = 10'h073;
        mem[20] = 10'h007;
        mem[21] = 10'h0bc;
        mem[22] = 10'h1bf;
        mem[23] = 10'h236;
        mem[24] = 10'h131;
        mem[25] = 10'h369;
        mem[26] = 10'h258;
        mem[27] = 10'h3bb;
        mem[28] = 10'h1cd;
        mem[29] = 10'h3a5;
        mem[30] = 10'h38a;
        mem[31] = 10'h1d5;
        mem[32] = 10'h3b9;
        mem[33] = 10'h1ad;
        mem[34] = 10'h0bb;
        mem[35] = 10'h2ae;
        mem[36] = 10'h3d6;
        mem[37] = 10'h359;
        mem[38] = 10'h302;
        mem[39] = 10'h34a;
        mem[40] = 10'h1c8;
        mem[41] = 10'h318;
        mem[42] = 10'h0b4;
        mem[43] = 10'h263;
        mem[44] = 10'h2f5;
        mem[45] = 10'h0c7;
        mem[46] = 10'h0a5;
        mem[47] = 10'h070;
        mem[48] = 10'h29e;
        mem[49] = 10'h3fd;
        mem[50] = 10'h2af;
        mem[51] = 10'h150;
        mem[52] = 10'h1ab;
        mem[53] = 10'h33b;
        mem[54] = 10'h24b;
        mem[55] = 10'h091;
        mem[56] = 10'h2a6;
        mem[57] = 10'h02d;
        mem[58] = 10'h32e;
        mem[59] = 10'h351;
        mem[60] = 10'h1dd;
        mem[61] = 10'h288;
        mem[62] = 10'h3d5;
        mem[63] = 10'h1c2;
        mem[64] = 10'h1a9;
        mem[65] = 10'h336;
        mem[66] = 10'h02f;
        mem[67] = 10'h02b;
        mem[68] = 10'h16a;
        mem[69] = 10'h21d;
        mem[70] = 10'h3f3;
        mem[71] = 10'h054;
        mem[72] = 10'h0b6;
        mem[73] = 10'h25d;
        mem[74] = 10'h3fe;
        mem[75] = 10'h246;
        mem[76] = 10'h134;
        mem[77] = 10'h3f2;
        mem[78] = 10'h055;
        mem[79] = 10'h09b;
        mem[80] = 10'h3bd;
        mem[81] = 10'h0c4;
        mem[82] = 10'h1de;
        mem[83] = 10'h170;
        mem[84] = 10'h034;
        mem[85] = 10'h321;
        mem[86] = 10'h162;
        mem[87] = 10'h3ba;
        mem[88] = 10'h1d8;
        mem[89] = 10'h3a1;
        mem[90] = 10'h2b0;
        mem[91] = 10'h2be;
        mem[92] = 10'h371;
        mem[93] = 10'h174;
        mem[94] = 10'h105;
        mem[95] = 10'h25f;
        mem[96] = 10'h0b1;
        mem[97] = 10'h2b9;
        mem[98] = 10'h2ca;
        mem[99] = 10'h32b;
        mem[100] = 10'h056;
        mem[101] = 10'h240;
        mem[102] = 10'h08f;
        mem[103] = 10'h193;
        mem[104] = 10'h192;
        mem[105] = 10'h340;
        mem[106] = 10'h182;
        mem[107] = 10'h2a7;
        mem[108] = 10'h2e1;
        mem[109] = 10'h0a2;
        mem[110] = 10'h04a;
        mem[111] = 10'h2bf;
        mem[112] = 10'h223;
        mem[113] = 10'h13c;
        mem[114] = 10'h275;
        mem[115] = 10'h32d;
        mem[116] = 10'h14e;
        mem[117] = 10'h1f2;
        mem[118] = 10'h358;
        mem[119] = 10'h18e;
        mem[120] = 10'h244;
        mem[121] = 10'h016;
        mem[122] = 10'h146;
        mem[123] = 10'h23e;
        mem[124] = 10'h285;
        mem[125] = 10'h2ea;
        mem[126] = 10'h0e6;
        mem[127] = 10'h19d;
        mem[128] = 10'h0f7;
        mem[129] = 10'h12f;
        mem[130] = 10'h305;
        mem[131] = 10'h15b;
        mem[132] = 10'h21c;
        mem[133] = 10'h3db;
        mem[134] = 10'h147;
        mem[135] = 10'h029;
        mem[136] = 10'h1fa;
        mem[137] = 10'h2d4;
        mem[138] = 10'h18f;
        mem[139] = 10'h2ad;
        mem[140] = 10'h230;
        mem[141] = 10'h327;
        mem[142] = 10'h383;
        mem[143] = 10'h206;
        mem[144] = 10'h391;
        mem[145] = 10'h179;
        mem[146] = 10'h18d;
        mem[147] = 10'h30e;
        mem[148] = 10'h19e;
        mem[149] = 10'h06b;
        mem[150] = 10'h0d1;
        mem[151] = 10'h108;
        mem[152] = 10'h104;
        mem[153] = 10'h0ab;
        mem[154] = 10'h110;
        mem[155] = 10'h20e;
        mem[156] = 10'h2ba;
        mem[157] = 10'h35e;
        mem[158] = 10'h37f;
        mem[159] = 10'h07c;
        mem[160] = 10'h265;
        mem[161] = 10'h07e;
        mem[162] = 10'h0f9;
        mem[163] = 10'h01c;
        mem[164] = 10'h26b;
        mem[165] = 10'h038;
        mem[166] = 10'h12b;
        mem[167] = 10'h200;
        mem[168] = 10'h3b1;
        mem[169] = 10'h16b;
        mem[170] = 10'h16c;
        mem[171] = 10'h07a;
        mem[172] = 10'h35f;
        mem[173] = 10'h1aa;
        mem[174] = 10'h2c4;
        mem[175] = 10'h119;
        mem[176] = 10'h3e1;
        mem[177] = 10'h178;
        mem[178] = 10'h069;
        mem[179] = 10'h02e;
        mem[180] = 10'h30d;
        mem[181] = 10'h009;
        mem[182] = 10'h2db;
        mem[183] = 10'h385;
        mem[184] = 10'h1e9;
        mem[185] = 10'h376;
        mem[186] = 10'h0c0;
        mem[187] = 10'h06f;
        mem[188] = 10'h3d0;
        mem[189] = 10'h3c8;
        mem[190] = 10'h163;
        mem[191] = 10'h388;
        mem[192] = 10'h0d6;
        mem[193] = 10'h323;
        mem[194] = 10'h2df;
        mem[195] = 10'h167;
        mem[196] = 10'h175;
        mem[197] = 10'h083;
        mem[198] = 10'h074;
        mem[199] = 10'h08b;
        mem[200] = 10'h11b;
        mem[201] = 10'h2f2;
        mem[202] = 10'h1f3;
        mem[203] = 10'h11a;
        mem[204] = 10'h2a5;
        mem[205] = 10'h24e;
        mem[206] = 10'h0c1;
        mem[207] = 10'h209;
        mem[208] = 10'h190;
        mem[209] = 10'h1d9;
        mem[210] = 10'h303;
        mem[211] = 10'h080;
        mem[212] = 10'h349;
        mem[213] = 10'h272;
        mem[214] = 10'h256;
        mem[215] = 10'h35a;
        mem[216] = 10'h082;
        mem[217] = 10'h3ea;
        mem[218] = 10'h149;
        mem[219] = 10'h28c;
        mem[220] = 10'h031;
        mem[221] = 10'h101;
        mem[222] = 10'h255;
        mem[223] = 10'h26c;
        mem[224] = 10'h26f;
        mem[225] = 10'h113;
        mem[226] = 10'h22d;
        mem[227] = 10'h36c;
        mem[228] = 10'h050;
        mem[229] = 10'h012;
        mem[230] = 10'h386;
        mem[231] = 10'h06e;
        mem[232] = 10'h027;
        mem[233] = 10'h291;
        mem[234] = 10'h34f;
        mem[235] = 10'h392;
        mem[236] = 10'h3ec;
        mem[237] = 10'h22b;
        mem[238] = 10'h23d;
        mem[239] = 10'h195;
        mem[240] = 10'h138;
        mem[241] = 10'h2b4;
        mem[242] = 10'h3b4;
        mem[243] = 10'h14c;
        mem[244] = 10'h2a1;
        mem[245] = 10'h09f;
        mem[246] = 10'h3e6;
        mem[247] = 10'h1e3;
        mem[248] = 10'h20b;
        mem[249] = 10'h023;
        mem[250] = 10'h0a1;
        mem[251] = 10'h2bb;
        mem[252] = 10'h38c;
        mem[253] = 10'h10e;
        mem[254] = 10'h13e;
        mem[255] = 10'h251;
        mem[256] = 10'h3cc;
        mem[257] = 10'h123;
        mem[258] = 10'h1fb;
        mem[259] = 10'h3d1;
        mem[260] = 10'h31d;
        mem[261] = 10'h29d;
        mem[262] = 10'h316;
        mem[263] = 10'h1d7;
        mem[264] = 10'h207;
        mem[265] = 10'h130;
        mem[266] = 10'h350;
        mem[267] = 10'h143;
        mem[268] = 10'h2b2;
        mem[269] = 10'h228;
        mem[270] = 10'h3c3;
        mem[271] = 10'h395;
        mem[272] = 10'h1ce;
        mem[273] = 10'h3f5;
        mem[274] = 10'h382;
        mem[275] = 10'h0db;
        mem[276] = 10'h10b;
        mem[277] = 10'h0fe;
        mem[278] = 10'h357;
        mem[279] = 10'h217;
        mem[280] = 10'h2f6;
        mem[281] = 10'h1d0;
        mem[282] = 10'h252;
        mem[283] = 10'h269;
        mem[284] = 10'h0bd;
        mem[285] = 10'h032;
        mem[286] = 10'h06d;
        mem[287] = 10'h24c;
        mem[288] = 10'h0e1;
        mem[289] = 10'h04e;
        mem[290] = 10'h354;
        mem[291] = 10'h36f;
        mem[292] = 10'h135;
        mem[293] = 10'h37e;
        mem[294] = 10'h3c4;
        mem[295] = 10'h237;
        mem[296] = 10'h21b;
        mem[297] = 10'h030;
        mem[298] = 10'h3da;
        mem[299] = 10'h0b0;
        mem[300] = 10'h144;
        mem[301] = 10'h14f;
        mem[302] = 10'h124;
        mem[303] = 10'h05e;
        mem[304] = 10'h211;
        mem[305] = 10'h374;
        mem[306] = 10'h384;
        mem[307] = 10'h099;
        mem[308] = 10'h037;
        mem[309] = 10'h3d9;
        mem[310] = 10'h0f3;
        mem[311] = 10'h2e8;
        mem[312] = 10'h15e;
        mem[313] = 10'h3bc;
        mem[314] = 10'h194;
        mem[315] = 10'h189;
        mem[316] = 10'h2cf;
        mem[317] = 10'h159;
        mem[318] = 10'h061;
        mem[319] = 10'h238;
        mem[320] = 10'h08a;
        mem[321] = 10'h087;
        mem[322] = 10'h267;
        mem[323] = 10'h18c;
        mem[324] = 10'h286;
        mem[325] = 10'h2dd;
        mem[326] = 10'h094;
        mem[327] = 10'h12a;
        mem[328] = 10'h341;
        mem[329] = 10'h1e2;
        mem[330] = 10'h249;
        mem[331] = 10'h346;
        mem[332] = 10'h1c4;
        mem[333] = 10'h365;
        mem[334] = 10'h052;
        mem[335] = 10'h096;
        mem[336] = 10'h3be;
        mem[337] = 10'h2c8;
        mem[338] = 10'h020;
        mem[339] = 10'h1be;
        mem[340] = 10'h026;
        mem[341] = 10'h0e5;
        mem[342] = 10'h3aa;
        mem[343] = 10'h1b3;
        mem[344] = 10'h3b7;
        mem[345] = 10'h245;
        mem[346] = 10'h27b;
        mem[347] = 10'h06a;
        mem[348] = 10'h30f;
        mem[349] = 10'h118;
        mem[350] = 10'h2d8;
        mem[351] = 10'h0ef;
        mem[352] = 10'h338;
        mem[353] = 10'h15c;
        mem[354] = 10'h2dc;
        mem[355] = 10'h320;
        mem[356] = 10'h3bf;
        mem[357] = 10'h2e6;
        mem[358] = 10'h16d;
        mem[359] = 10'h37a;
        mem[360] = 10'h01a;
        mem[361] = 10'h33f;
        mem[362] = 10'h043;
        mem[363] = 10'h107;
        mem[364] = 10'h2e0;
        mem[365] = 10'h35c;
        mem[366] = 10'h3cd;
        mem[367] = 10'h39c;
        mem[368] = 10'h0ff;
        mem[369] = 10'h156;
        mem[370] = 10'h0f2;
        mem[371] = 10'h18b;
        mem[372] = 10'h126;
        mem[373] = 10'h242;
        mem[374] = 10'h0e4;
        mem[375] = 10'h045;
        mem[376] = 10'h2f3;
        mem[377] = 10'h30b;
        mem[378] = 10'h283;
        mem[379] = 10'h025;
        mem[380] = 10'h039;
        mem[381] = 10'h17f;
        mem[382] = 10'h25e;
        mem[383] = 10'h2bc;
        mem[384] = 10'h198;
        mem[385] = 10'h2ff;
        mem[386] = 10'h281;
        mem[387] = 10'h0fd;
        mem[388] = 10'h3e8;
        mem[389] = 10'h229;
        mem[390] = 10'h04d;
        mem[391] = 10'h2b1;
        mem[392] = 10'h3ad;
        mem[393] = 10'h03e;
        mem[394] = 10'h1ac;
        mem[395] = 10'h25a;
        mem[396] = 10'h362;
        mem[397] = 10'h0cb;
        mem[398] = 10'h010;
        mem[399] = 10'h312;
        mem[400] = 10'h333;
        mem[401] = 10'h3a7;
        mem[402] = 10'h014;
        mem[403] = 10'h003;
        mem[404] = 10'h247;
        mem[405] = 10'h271;
        mem[406] = 10'h157;
        mem[407] = 10'h2b6;
        mem[408] = 10'h1b8;
        mem[409] = 10'h231;
        mem[410] = 10'h243;
        mem[411] = 10'h3de;
        mem[412] = 10'h287;
        mem[413] = 10'h3d4;
        mem[414] = 10'h202;
        mem[415] = 10'h0a4;
        mem[416] = 10'h0f6;
        mem[417] = 10'h334;
        mem[418] = 10'h0b8;
        mem[419] = 10'h1af;
        mem[420] = 10'h364;
        mem[421] = 10'h121;
        mem[422] = 10'h3f6;
        mem[423] = 10'h2c3;
        mem[424] = 10'h0fc;
        mem[425] = 10'h197;
        mem[426] = 10'h2d0;
        mem[427] = 10'h3b5;
        mem[428] = 10'h2ec;
        mem[429] = 10'h3c6;
        mem[430] = 10'h11c;
        mem[431] = 10'h0b9;
        mem[432] = 10'h19a;
        mem[433] = 10'h148;
        mem[434] = 10'h2cb;
        mem[435] = 10'h373;
        mem[436] = 10'h31a;
        mem[437] = 10'h38d;
        mem[438] = 10'h19b;
        mem[439] = 10'h345;
        mem[440] = 10'h394;
        mem[441] = 10'h018;
        mem[442] = 10'h0eb;
        mem[443] = 10'h3a4;
        mem[444] = 10'h279;
        mem[445] = 10'h356;
        mem[446] = 10'h2fb;
        mem[447] = 10'h2cd;
        mem[448] = 10'h22c;
        mem[449] = 10'h114;
        mem[450] = 10'h266;
        mem[451] = 10'h220;
        mem[452] = 10'h21f;
        mem[453] = 10'h115;
        mem[454] = 10'h186;
        mem[455] = 10'h076;
        mem[456] = 10'h304;
        mem[457] = 10'h0a6;
        mem[458] = 10'h3ac;
        mem[459] = 10'h01b;
        mem[460] = 10'h3f7;
        mem[461] = 10'h2d1;
        mem[462] = 10'h0c5;
        mem[463] = 10'h370;
        mem[464] = 10'h307;
        mem[465] = 10'h053;
        mem[466] = 10'h29c;
        mem[467] = 10'h284;
        mem[468] = 10'h2aa;
        mem[469] = 10'h03d;
        mem[470] = 10'h20f;
        mem[471] = 10'h28e;
        mem[472] = 10'h199;
        mem[473] = 10'h23c;
        mem[474] = 10'h27c;
        mem[475] = 10'h0d2;
        mem[476] = 10'h222;
        mem[477] = 10'h1e1;
        mem[478] = 10'h31f;
        mem[479] = 10'h280;
        mem[480] = 10'h05f;
        mem[481] = 10'h13f;
        mem[482] = 10'h1bb;
        mem[483] = 10'h1a1;
        mem[484] = 10'h00d;
        mem[485] = 10'h33a;
        mem[486] = 10'h344;
        mem[487] = 10'h1ed;
        mem[488] = 10'h2e5;
        mem[489] = 10'h381;
        mem[490] = 10'h05a;
        mem[491] = 10'h1cb;
        mem[492] = 10'h139;
        mem[493] = 10'h397;
        mem[494] = 10'h04c;
        mem[495] = 10'h075;
        mem[496] = 10'h152;
        mem[497] = 10'h2e3;
        mem[498] = 10'h3c5;
        mem[499] = 10'h01e;
        mem[500] = 10'h173;
        mem[501] = 10'h0d9;
        mem[502] = 10'h2c1;
        mem[503] = 10'h268;
        mem[504] = 10'h2c7;
        mem[505] = 10'h187;
        mem[506] = 10'h2c6;
        mem[507] = 10'h2a3;
        mem[508] = 10'h1d2;
        mem[509] = 10'h23b;
        mem[510] = 10'h319;
        mem[511] = 10'h298;
        mem[512] = 10'h127;
        mem[513] = 10'h1bc;
        mem[514] = 10'h081;
        mem[515] = 10'h044;
        mem[516] = 10'h214;
        mem[517] = 10'h32a;
        mem[518] = 10'h028;
        mem[519] = 10'h142;
        mem[520] = 10'h23a;
        mem[521] = 10'h060;
        mem[522] = 10'h250;
        mem[523] = 10'h111;
        mem[524] = 10'h117;
        mem[525] = 10'h02a;
        mem[526] = 10'h353;
        mem[527] = 10'h38f;
        mem[528] = 10'h315;
        mem[529] = 10'h0a8;
        mem[530] = 10'h0cf;
        mem[531] = 10'h3fc;
        mem[532] = 10'h262;
        mem[533] = 10'h3f9;
        mem[534] = 10'h232;
        mem[535] = 10'h006;
        mem[536] = 10'h25c;
        mem[537] = 10'h0c2;
        mem[538] = 10'h2a2;
        mem[539] = 10'h30c;
        mem[540] = 10'h2b5;
        mem[541] = 10'h261;
        mem[542] = 10'h0d7;
        mem[543] = 10'h0cd;
        mem[544] = 10'h313;
        mem[545] = 10'h26e;
        mem[546] = 10'h128;
        mem[547] = 10'h093;
        mem[548] = 10'h39e;
        mem[549] = 10'h3f1;
        mem[550] = 10'h3a2;
        mem[551] = 10'h3dc;
        mem[552] = 10'h1b0;
        mem[553] = 10'h2a9;
        mem[554] = 10'h1ef;
        mem[555] = 10'h0e0;
        mem[556] = 10'h2e2;
        mem[557] = 10'h180;
        mem[558] = 10'h1ba;
        mem[559] = 10'h0ae;
        mem[560] = 10'h37b;
        mem[561] = 10'h39b;
        mem[562] = 10'h1b1;
        mem[563] = 10'h01f;
        mem[564] = 10'h330;
        mem[565] = 10'h3c0;
        mem[566] = 10'h29b;
        mem[567] = 10'h078;
        mem[568] = 10'h3b8;
        mem[569] = 10'h161;
        mem[570] = 10'h290;
        mem[571] = 10'h295;
        mem[572] = 10'h097;
        mem[573] = 10'h3ca;
        mem[574] = 10'h377;
        mem[575] = 10'h13d;
        mem[576] = 10'h3ef;
        mem[577] = 10'h0f4;
        mem[578] = 10'h270;
        mem[579] = 10'h38e;
        mem[580] = 10'h09c;
        mem[581] = 10'h3e5;
        mem[582] = 10'h2d3;
        mem[583] = 10'h0d4;
        mem[584] = 10'h322;
        mem[585] = 10'h116;
        mem[586] = 10'h1f1;
        mem[587] = 10'h342;
        mem[588] = 10'h019;
        mem[589] = 10'h219;
        mem[590] = 10'h0cc;
        mem[591] = 10'h248;
        mem[592] = 10'h1cf;
        mem[593] = 10'h160;
        mem[594] = 10'h3b0;
        mem[595] = 10'h068;
        mem[596] = 10'h2fd;
        mem[597] = 10'h294;
        mem[598] = 10'h264;
        mem[599] = 10'h2d5;
        mem[600] = 10'h122;
        mem[601] = 10'h0be;
        mem[602] = 10'h16f;
        mem[603] = 10'h1ec;
        mem[604] = 10'h29f;
        mem[605] = 10'h17e;
        mem[606] = 10'h2de;
        mem[607] = 10'h015;
        mem[608] = 10'h39f;
        mem[609] = 10'h208;
        mem[610] = 10'h2f4;
        mem[611] = 10'h0fa;
        mem[612] = 10'h0f5;
        mem[613] = 10'h337;
        mem[614] = 10'h10a;
        mem[615] = 10'h28b;
        mem[616] = 10'h085;
        mem[617] = 10'h299;
        mem[618] = 10'h22a;
        mem[619] = 10'h0a0;
        mem[620] = 10'h225;
        mem[621] = 10'h29a;
        mem[622] = 10'h1fd;
        mem[623] = 10'h1da;
        mem[624] = 10'h2e7;
        mem[625] = 10'h1ae;
        mem[626] = 10'h0e9;
        mem[627] = 10'h218;
        mem[628] = 10'h254;
        mem[629] = 10'h0ad;
        mem[630] = 10'h11d;
        mem[631] = 10'h01d;
        mem[632] = 10'h1e0;
        mem[633] = 10'h1a4;
        mem[634] = 10'h2c5;
        mem[635] = 10'h2ed;
        mem[636] = 10'h31e;
        mem[637] = 10'h03a;
        mem[638] = 10'h3c2;
        mem[639] = 10'h3fb;
        mem[640] = 10'h0dd;
        mem[641] = 10'h2a4;
        mem[642] = 10'h15a;
        mem[643] = 10'h15f;
        mem[644] = 10'h3e7;
        mem[645] = 10'h1bd;
        mem[646] = 10'h067;
        mem[647] = 10'h1a3;
        mem[648] = 10'h1d4;
        mem[649] = 10'h0bf;
        mem[650] = 10'h331;
        mem[651] = 10'h311;
        mem[652] = 10'h339;
        mem[653] = 10'h011;
        mem[654] = 10'h224;
        mem[655] = 10'h0b2;
        mem[656] = 10'h0da;
        mem[657] = 10'h1fe;
        mem[658] = 10'h276;
        mem[659] = 10'h1b7;
        mem[660] = 10'h095;
        mem[661] = 10'h0f8;
        mem[662] = 10'h293;
        mem[663] = 10'h2ab;
        mem[664] = 10'h2d6;
        mem[665] = 10'h0e8;
        mem[666] = 10'h39d;
        mem[667] = 10'h2a8;
        mem[668] = 10'h1c7;
        mem[669] = 10'h289;
        mem[670] = 10'h086;
        mem[671] = 10'h00b;
        mem[672] = 10'h28d;
        mem[673] = 10'h2e4;
        mem[674] = 10'h106;
        mem[675] = 10'h0ea;
        mem[676] = 10'h04b;
        mem[677] = 10'h05b;
        mem[678] = 10'h3fa;
        mem[679] = 10'h0b7;
        mem[680] = 10'h3a0;
        mem[681] = 10'h3c9;
        mem[682] = 10'h3eb;
        mem[683] = 10'h239;
        mem[684] = 10'h23f;
        mem[685] = 10'h0d8;
        mem[686] = 10'h277;
        mem[687] = 10'h177;
        mem[688] = 10'h2c9;
        mem[689] = 10'h36b;
        mem[690] = 10'h0ca;
        mem[691] = 10'h00e;
        mem[692] = 10'h387;
        mem[693] = 10'h102;
        mem[694] = 10'h136;
        mem[695] = 10'h3e3;
        mem[696] = 10'h35b;
        mem[697] = 10'h059;
        mem[698] = 10'h278;
        mem[699] = 10'h2eb;
        mem[700] = 10'h30a;
        mem[701] = 10'h2ef;
        mem[702] = 10'h1f5;
        mem[703] = 10'h1d6;
        mem[704] = 10'h308;
        mem[705] = 10'h10c;
        mem[706] = 10'h2fa;
        mem[707] = 10'h09e;
        mem[708] = 10'h2d7;
        mem[709] = 10'h31c;
        mem[710] = 10'h1c1;
        mem[711] = 10'h06c;
        mem[712] = 10'h2fc;
        mem[713] = 10'h375;
        mem[714] = 10'h0ec;
        mem[715] = 10'h301;
        mem[716] = 10'h393;
        mem[717] = 10'h36e;
        mem[718] = 10'h066;
        mem[719] = 10'h20a;
        mem[720] = 10'h005;
        mem[721] = 10'h2d2;
        mem[722] = 10'h041;
        mem[723] = 10'h188;
        mem[724] = 10'h274;
        mem[725] = 10'h022;
        mem[726] = 10'h141;
        mem[727] = 10'h098;
        mem[728] = 10'h257;
        mem[729] = 10'h3e4;
        mem[730] = 10'h17a;
        mem[731] = 10'h3cf;
        mem[732] = 10'h28a;
        mem[733] = 10'h0e2;
        mem[734] = 10'h324;
        mem[735] = 10'h0ee;
        mem[736] = 10'h1f0;
        mem[737] = 10'h216;
        mem[738] = 10'h17d;
        mem[739] = 10'h02c;
        mem[740] = 10'h201;
        mem[741] = 10'h0df;
        mem[742] = 10'h1fc;
        mem[743] = 10'h0a9;
        mem[744] = 10'h017;
        mem[745] = 10'h03f;
        mem[746] = 10'h3d3;
        mem[747] = 10'h103;
        mem[748] = 10'h11e;
        mem[749] = 10'h3d2;
        mem[750] = 10'h259;
        mem[751] = 10'h063;
        mem[752] = 10'h205;
        mem[753] = 10'h25b;
        mem[754] = 10'h04f;
        mem[755] = 10'h24a;
        mem[756] = 10'h14a;
        mem[757] = 10'h3cb;
        mem[758] = 10'h1a7;
        mem[759] = 10'h0c9;
        mem[760] = 10'h27f;
        mem[761] = 10'h1a8;
        mem[762] = 10'h0b3;
        mem[763] = 10'h089;
        mem[764] = 10'h3e2;
        mem[765] = 10'h241;
        mem[766] = 10'h2b7;
        mem[767] = 10'h051;
        mem[768] = 10'h035;
        mem[769] = 10'h0e7;
        mem[770] = 10'h1b4;
        mem[771] = 10'h12c;
        mem[772] = 10'h191;
        mem[773] = 10'h347;
        mem[774] = 10'h008;
        mem[775] = 10'h366;
        mem[776] = 10'h092;
        mem[777] = 10'h3ce;
        mem[778] = 10'h08c;
        mem[779] = 10'h21a;
        mem[780] = 10'h28f;
        mem[781] = 10'h348;
        mem[782] = 10'h09d;
        mem[783] = 10'h05c;
        mem[784] = 10'h389;
        mem[785] = 10'h36a;
        mem[786] = 10'h22e;
        mem[787] = 10'h140;
        mem[788] = 10'h378;
        mem[789] = 10'h3ab;
        mem[790] = 10'h32f;
        mem[791] = 10'h07d;
        mem[792] = 10'h181;
        mem[793] = 10'h0f0;
        mem[794] = 10'h2d9;
        mem[795] = 10'h260;
        mem[796] = 10'h1a5;
        mem[797] = 10'h227;
        mem[798] = 10'h3df;
        mem[799] = 10'h27a;
        mem[800] = 10'h3a3;
        mem[801] = 10'h196;
        mem[802] = 10'h26d;
        mem[803] = 10'h151;
        mem[804] = 10'h3ae;
        mem[805] = 10'h0c3;
        mem[806] = 10'h363;
        mem[807] = 10'h1ca;
        mem[808] = 10'h398;
        mem[809] = 10'h352;
        mem[810] = 10'h27e;
        mem[811] = 10'h004;
        mem[812] = 10'h154;
        mem[813] = 10'h1b9;
        mem[814] = 10'h13a;
        mem[815] = 10'h049;
        mem[816] = 10'h013;
        mem[817] = 10'h11f;
        mem[818] = 10'h37c;
        mem[819] = 10'h0ba;
        mem[820] = 10'h27d;
        mem[821] = 10'h024;
        mem[822] = 10'h184;
        mem[823] = 10'h34c;
        mem[824] = 10'h1f7;
        mem[825] = 10'h155;
        mem[826] = 10'h048;
        mem[827] = 10'h166;
        mem[828] = 10'h15d;
        mem[829] = 10'h19c;
        mem[830] = 10'h0e3;
        mem[831] = 10'h19f;
        mem[832] = 10'h396;
        mem[833] = 10'h335;
        mem[834] = 10'h1a6;
        mem[835] = 10'h1ff;
        mem[836] = 10'h0aa;
        mem[837] = 10'h204;
        mem[838] = 10'h10d;
        mem[839] = 10'h00c;
        mem[840] = 10'h292;
        mem[841] = 10'h328;
        mem[842] = 10'h39a;
        mem[843] = 10'h0ac;
        mem[844] = 10'h1c3;
        mem[845] = 10'h399;
        mem[846] = 10'h3a6;
        mem[847] = 10'h213;
        mem[848] = 10'h1cc;
        mem[849] = 10'h35d;
        mem[850] = 10'h03c;
        mem[851] = 10'h17c;
        mem[852] = 10'h1a0;
        mem[853] = 10'h1df;
        mem[854] = 10'h002;
        mem[855] = 10'h1a2;
        mem[856] = 10'h3a9;
        mem[857] = 10'h235;
        mem[858] = 10'h14d;
        mem[859] = 10'h3d7;
        mem[860] = 10'h24f;
        mem[861] = 10'h37d;
        mem[862] = 10'h210;
        mem[863] = 10'h2f8;
        mem[864] = 10'h001;
        mem[865] = 10'h367;
        mem[866] = 10'h10f;
        mem[867] = 10'h2f1;
        mem[868] = 10'h2cc;
        mem[869] = 10'h0fb;
        mem[870] = 10'h226;
        mem[871] = 10'h0a7;
        mem[872] = 10'h176;
        mem[873] = 10'h1c6;
        mem[874] = 10'h2bd;
        mem[875] = 10'h3b2;
        mem[876] = 10'h047;
        mem[877] = 10'h0b5;
        mem[878] = 10'h343;
        mem[879] = 10'h1f6;
        mem[880] = 10'h253;
        mem[881] = 10'h203;
        mem[882] = 10'h14b;
        mem[883] = 10'h3ed;
        mem[884] = 10'h1e5;
        mem[885] = 10'h129;
        mem[886] = 10'h065;
        mem[887] = 10'h212;
        mem[888] = 10'h1eb;
        mem[889] = 10'h31b;
        mem[890] = 10'h0f1;
        mem[891] = 10'h361;
        mem[892] = 10'h2c0;
        mem[893] = 10'h133;
        mem[894] = 10'h0d0;
        mem[895] = 10'h071;
        mem[896] = 10'h168;
        mem[897] = 10'h1d1;
        mem[898] = 10'h036;
        mem[899] = 10'h2ce;
        mem[900] = 10'h215;
        mem[901] = 10'h1f4;
        mem[902] = 10'h0ce;
        mem[903] = 10'h1c0;
        mem[904] = 10'h1c5;
        mem[905] = 10'h32c;
        mem[906] = 10'h3f4;
        mem[907] = 10'h296;
        mem[908] = 10'h2da;
        mem[909] = 10'h062;
        mem[910] = 10'h3ee;
        mem[911] = 10'h390;
        mem[912] = 10'h171;
        mem[913] = 10'h0ed;
        mem[914] = 10'h20c;
        mem[915] = 10'h079;
        mem[916] = 10'h040;
        mem[917] = 10'h169;
        mem[918] = 10'h03b;
        mem[919] = 10'h021;
        mem[920] = 10'h3e0;
        mem[921] = 10'h2f7;
        mem[922] = 10'h2fe;
        mem[923] = 10'h22f;
        mem[924] = 10'h1d3;
        mem[925] = 10'h05d;
        mem[926] = 10'h1f9;
        mem[927] = 10'h0af;
        mem[928] = 10'h3ff;
        mem[929] = 10'h38b;
        mem[930] = 10'h0de;
        mem[931] = 10'h09a;
        mem[932] = 10'h300;
        mem[933] = 10'h24d;
        mem[934] = 10'h233;
        mem[935] = 10'h153;
        mem[936] = 10'h1b5;
        mem[937] = 10'h221;
        mem[938] = 10'h2ee;
        mem[939] = 10'h0a3;
        mem[940] = 10'h234;
        mem[941] = 10'h368;
        mem[942] = 10'h2f9;
        mem[943] = 10'h33d;
        mem[944] = 10'h326;
        mem[945] = 10'h282;
        mem[946] = 10'h1b6;
        mem[947] = 10'h3f8;
        mem[948] = 10'h317;
        mem[949] = 10'h3f0;
        mem[950] = 10'h36d;
        mem[951] = 10'h273;
        mem[952] = 10'h3af;
        mem[953] = 10'h137;
        mem[954] = 10'h3d8;
        mem[955] = 10'h3c1;
        mem[956] = 10'h17b;
        mem[957] = 10'h08e;
        mem[958] = 10'h064;
        mem[959] = 10'h183;
        mem[960] = 10'h297;
        mem[961] = 10'h2a0;
        mem[962] = 10'h380;
        mem[963] = 10'h057;
        mem[964] = 10'h158;
        mem[965] = 10'h1f8;
        mem[966] = 10'h2b3;
        mem[967] = 10'h00f;
        mem[968] = 10'h34b;
        mem[969] = 10'h2f0;
        mem[970] = 10'h33c;
        mem[971] = 10'h314;
        mem[972] = 10'h172;
        mem[973] = 10'h185;
        mem[974] = 10'h2ac;
        mem[975] = 10'h120;
        mem[976] = 10'h088;
        mem[977] = 10'h0d5;
        mem[978] = 10'h164;
        mem[979] = 10'h058;
        mem[980] = 10'h0d3;
        mem[981] = 10'h3e9;
        mem[982] = 10'h20d;
        mem[983] = 10'h1ee;
        mem[984] = 10'h109;
        mem[985] = 10'h332;
        mem[986] = 10'h34d;
        mem[987] = 10'h13b;
        mem[988] = 10'h145;
        mem[989] = 10'h309;
        mem[990] = 10'h072;
        mem[991] = 10'h3dd;
        mem[992] = 10'h18a;
        mem[993] = 10'h355;
        mem[994] = 10'h0c6;
        mem[995] = 10'h1e4;
        mem[996] = 10'h1b2;
        mem[997] = 10'h125;
        mem[998] = 10'h3b6;
        mem[999] = 10'h084;
        mem[1000] = 10'h1db;
        mem[1001] = 10'h000;
        mem[1002] = 10'h2b8;
        mem[1003] = 10'h0c8;
        mem[1004] = 10'h077;
        mem[1005] = 10'h33e;
        mem[1006] = 10'h08d;
        mem[1007] = 10'h12e;
        mem[1008] = 10'h3b3;
        mem[1009] = 10'h100;
        mem[1010] = 10'h090;
        mem[1011] = 10'h3c7;
        mem[1012] = 10'h26a;
        mem[1013] = 10'h112;
        mem[1014] = 10'h2c2;
        mem[1015] = 10'h12d;
        mem[1016] = 10'h1e8;
        mem[1017] = 10'h033;
        mem[1018] = 10'h310;
        mem[1019] = 10'h2e9;
        mem[1020] = 10'h360;
        mem[1021] = 10'h046;
        mem[1022] = 10'h165;
        mem[1023] = 10'h1e7;
    end
endmodule

module odo_sbox_large2(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    (* ram_style = "block" *) reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h278;
        mem[1] = 10'h17e;
        mem[2] = 10'h348;
        mem[3] = 10'h168;
        mem[4] = 10'h1f4;
        mem[5] = 10'h367;
        mem[6] = 10'h016;
        mem[7] = 10'h0ff;
        mem[8] = 10'h3f6;
        mem[9] = 10'h375;
        mem[10] = 10'h39e;
        mem[11] = 10'h250;
        mem[12] = 10'h1d4;
        mem[13] = 10'h319;
        mem[14] = 10'h114;
        mem[15] = 10'h3e1;
        mem[16] = 10'h18e;
        mem[17] = 10'h276;
        mem[18] = 10'h360;
        mem[19] = 10'h24e;
        mem[20] = 10'h248;
        mem[21] = 10'h103;
        mem[22] = 10'h2f9;
        mem[23] = 10'h0f7;
        mem[24] = 10'h142;
        mem[25] = 10'h09a;
        mem[26] = 10'h1ed;
        mem[27] = 10'h017;
        mem[28] = 10'h2cf;
        mem[29] = 10'h2e9;
        mem[30] = 10'h1c2;
        mem[31] = 10'h25d;
        mem[32] = 10'h140;
        mem[33] = 10'h10f;
        mem[34] = 10'h361;
        mem[35] = 10'h0f1;
        mem[36] = 10'h1a8;
        mem[37] = 10'h2aa;
        mem[38] = 10'h396;
        mem[39] = 10'h024;
        mem[40] = 10'h078;
        mem[41] = 10'h032;
        mem[42] = 10'h26f;
        mem[43] = 10'h138;
        mem[44] = 10'h306;
        mem[45] = 10'h230;
        mem[46] = 10'h193;
        mem[47] = 10'h08e;
        mem[48] = 10'h363;
        mem[49] = 10'h0f5;
        mem[50] = 10'h298;
        mem[51] = 10'h2bb;
        mem[52] = 10'h1b8;
        mem[53] = 10'h06d;
        mem[54] = 10'h3d9;
        mem[55] = 10'h350;
        mem[56] = 10'h10b;
        mem[57] = 10'h26b;
        mem[58] = 10'h112;
        mem[59] = 10'h3dd;
        mem[60] = 10'h000;
        mem[61] = 10'h0fe;
        mem[62] = 10'h272;
        mem[63] = 10'h2d6;
        mem[64] = 10'h356;
        mem[65] = 10'h013;
        mem[66] = 10'h3c2;
        mem[67] = 10'h172;
        mem[68] = 10'h159;
        mem[69] = 10'h23c;
        mem[70] = 10'h1f0;
        mem[71] = 10'h35e;
        mem[72] = 10'h058;
        mem[73] = 10'h13d;
        mem[74] = 10'h16b;
        mem[75] = 10'h2bf;
        mem[76] = 10'h376;
        mem[77] = 10'h150;
        mem[78] = 10'h1b0;
        mem[79] = 10'h12d;
        mem[80] = 10'h0c1;
        mem[81] = 10'h045;
        mem[82] = 10'h371;
        mem[83] = 10'h3a4;
        mem[84] = 10'h2b3;
        mem[85] = 10'h2c9;
        mem[86] = 10'h3a5;
        mem[87] = 10'h31f;
        mem[88] = 10'h01f;
        mem[89] = 10'h0e0;
        mem[90] = 10'h255;
        mem[91] = 10'h36d;
        mem[92] = 10'h006;
        mem[93] = 10'h3f0;
        mem[94] = 10'h2f2;
        mem[95] = 10'h1a2;
        mem[96] = 10'h1a6;
        mem[97] = 10'h143;
        mem[98] = 10'h008;
        mem[99] = 10'h183;
        mem[100] = 10'h2ad;
        mem[101] = 10'h11b;
        mem[102] = 10'h18f;
        mem[103] = 10'h0ae;
        mem[104] = 10'h352;
        mem[105] = 10'h1ab;
        mem[106] = 10'h3b4;
        mem[107] = 10'h2b9;
        mem[108] = 10'h1f5;
        mem[109] = 10'h2ed;
        mem[110] = 10'h038;
        mem[111] = 10'h266;
        mem[112] = 10'h0a0;
        mem[113] = 10'h20f;
        mem[114] = 10'h1a3;
        mem[115] = 10'h061;
        mem[116] = 10'h3b1;
        mem[117] = 10'h3d5;
        mem[118] = 10'h125;
        mem[119] = 10'h0a8;
        mem[120] = 10'h16c;
        mem[121] = 10'h246;
        mem[122] = 10'h232;
        mem[123] = 10'h001;
        mem[124] = 10'h0ce;
        mem[125] = 10'h06a;
        mem[126] = 10'h155;
        mem[127] = 10'h21e;
        mem[128] = 10'h054;
        mem[129] = 10'h02b;
        mem[130] = 10'h3b3;
        mem[131] = 10'h3c4;
        mem[132] = 10'h01c;
        mem[133] = 10'h294;
        mem[134] = 10'h33a;
        mem[135] = 10'h2a2;
        mem[136] = 10'h277;
        mem[137] = 10'h264;
        mem[138] = 10'h027;
        mem[139] = 10'h3c7;
        mem[140] = 10'h3cd;
        mem[141] = 10'h347;
        mem[142] = 10'h215;
        mem[143] = 10'h07d;
        mem[144] = 10'h313;
        mem[145] = 10'h39f;
        mem[146] = 10'h0ac;
        mem[147] = 10'h249;
        mem[148] = 10'h124;
        mem[149] = 10'h206;
        mem[150] = 10'h1c1;
        mem[151] = 10'h366;
        mem[152] = 10'h3de;
        mem[153] = 10'h34d;
        mem[154] = 10'h192;
        mem[155] = 10'h3d8;
        mem[156] = 10'h273;
        mem[157] = 10'h186;
        mem[158] = 10'h339;
        mem[159] = 10'h389;
        mem[160] = 10'h2c1;
        mem[161] = 10'h260;
        mem[162] = 10'h02e;
        mem[163] = 10'h32f;
        mem[164] = 10'h17a;
        mem[165] = 10'h329;
        mem[166] = 10'h145;
        mem[167] = 10'h27c;
        mem[168] = 10'h0d6;
        mem[169] = 10'h173;
        mem[170] = 10'h003;
        mem[171] = 10'h210;
        mem[172] = 10'h0af;
        mem[173] = 10'h20e;
        mem[174] = 10'h189;
        mem[175] = 10'h044;
        mem[176] = 10'h0a9;
        mem[177] = 10'h1b2;
        mem[178] = 10'h07e;
        mem[179] = 10'h3f5;
        mem[180] = 10'h207;
        mem[181] = 10'h27b;
        mem[182] = 10'h29e;
        mem[183] = 10'h086;
        mem[184] = 10'h0c4;
        mem[185] = 10'h2a0;
        mem[186] = 10'h072;
        mem[187] = 10'h34c;
        mem[188] = 10'h171;
        mem[189] = 10'h2ba;
        mem[190] = 10'h15e;
        mem[191] = 10'h146;
        mem[192] = 10'h1ba;
        mem[193] = 10'h1d8;
        mem[194] = 10'h383;
        mem[195] = 10'h213;
        mem[196] = 10'h3f8;
        mem[197] = 10'h285;
        mem[198] = 10'h0c6;
        mem[199] = 10'h228;
        mem[200] = 10'h237;
        mem[201] = 10'h0d2;
        mem[202] = 10'h0b5;
        mem[203] = 10'h00d;
        mem[204] = 10'h38f;
        mem[205] = 10'h0a4;
        mem[206] = 10'h0a3;
        mem[207] = 10'h0f3;
        mem[208] = 10'h162;
        mem[209] = 10'h205;
        mem[210] = 10'h25a;
        mem[211] = 10'h118;
        mem[212] = 10'h28e;
        mem[213] = 10'h15a;
        mem[214] = 10'h079;
        mem[215] = 10'h1ff;
        mem[216] = 10'h007;
        mem[217] = 10'h1a1;
        mem[218] = 10'h2f5;
        mem[219] = 10'h28f;
        mem[220] = 10'h1af;
        mem[221] = 10'h071;
        mem[222] = 10'h0cd;
        mem[223] = 10'h1fe;
        mem[224] = 10'h314;
        mem[225] = 10'h3d1;
        mem[226] = 10'h1c6;
        mem[227] = 10'h3fc;
        mem[228] = 10'h2d4;
        mem[229] = 10'h1b6;
        mem[230] = 10'h22f;
        mem[231] = 10'h34e;
        mem[232] = 10'h2ee;
        mem[233] = 10'h05b;
        mem[234] = 10'h020;
        mem[235] = 10'h0c7;
        mem[236] = 10'h093;
        mem[237] = 10'h084;
        mem[238] = 10'h07a;
        mem[239] = 10'h3a1;
        mem[240] = 10'h318;
        mem[241] = 10'h18a;
        mem[242] = 10'h057;
        mem[243] = 10'h3bd;
        mem[244] = 10'h065;
        mem[245] = 10'h323;
        mem[246] = 10'h369;
        mem[247] = 10'h381;
        mem[248] = 10'h316;
        mem[249] = 10'h060;
        mem[250] = 10'h187;
        mem[251] = 10'h048;
        mem[252] = 10'h342;
        mem[253] = 10'h297;
        mem[254] = 10'h3af;
        mem[255] = 10'h334;
        mem[256] = 10'h11e;
        mem[257] = 10'h201;
        mem[258] = 10'h00a;
        mem[259] = 10'h3c6;
        mem[260] = 10'h3be;
        mem[261] = 10'h01d;
        mem[262] = 10'h009;
        mem[263] = 10'h053;
        mem[264] = 10'h301;
        mem[265] = 10'h3a6;
        mem[266] = 10'h179;
        mem[267] = 10'h357;
        mem[268] = 10'h35d;
        mem[269] = 10'h094;
        mem[270] = 10'h31a;
        mem[271] = 10'h0f4;
        mem[272] = 10'h2bd;
        mem[273] = 10'h241;
        mem[274] = 10'h1de;
        mem[275] = 10'h19b;
        mem[276] = 10'h3d6;
        mem[277] = 10'h1d6;
        mem[278] = 10'h239;
        mem[279] = 10'h14b;
        mem[280] = 10'h0b7;
        mem[281] = 10'h300;
        mem[282] = 10'h174;
        mem[283] = 10'h10c;
        mem[284] = 10'h337;
        mem[285] = 10'h158;
        mem[286] = 10'h36e;
        mem[287] = 10'h2cc;
        mem[288] = 10'h131;
        mem[289] = 10'h119;
        mem[290] = 10'h128;
        mem[291] = 10'h267;
        mem[292] = 10'h039;
        mem[293] = 10'h11c;
        mem[294] = 10'h220;
        mem[295] = 10'h07c;
        mem[296] = 10'h19d;
        mem[297] = 10'h2d7;
        mem[298] = 10'h2de;
        mem[299] = 10'h33e;
        mem[300] = 10'h157;
        mem[301] = 10'h2e2;
        mem[302] = 10'h0b9;
        mem[303] = 10'h217;
        mem[304] = 10'h08d;
        mem[305] = 10'h3ac;
        mem[306] = 10'h021;
        mem[307] = 10'h0e6;
        mem[308] = 10'h176;
        mem[309] = 10'h1e2;
        mem[310] = 10'h268;
        mem[311] = 10'h333;
        mem[312] = 10'h324;
        mem[313] = 10'h26d;
        mem[314] = 10'h3e5;
        mem[315] = 10'h184;
        mem[316] = 10'h2e0;
        mem[317] = 10'h3ab;
        mem[318] = 10'h251;
        mem[319] = 10'h328;
        mem[320] = 10'h20c;
        mem[321] = 10'h1fc;
        mem[322] = 10'h27e;
        mem[323] = 10'h305;
        mem[324] = 10'h2da;
        mem[325] = 10'h00b;
        mem[326] = 10'h24f;
        mem[327] = 10'h351;
        mem[328] = 10'h0d3;
        mem[329] = 10'h132;
        mem[330] = 10'h359;
        mem[331] = 10'h37d;
        mem[332] = 10'h014;
        mem[333] = 10'h0b4;
        mem[334] = 10'h37e;
        mem[335] = 10'h0a5;
        mem[336] = 10'h099;
        mem[337] = 10'h108;
        mem[338] = 10'h1a4;
        mem[339] = 10'h136;
        mem[340] = 10'h098;
        mem[341] = 10'h393;
        mem[342] = 10'h144;
        mem[343] = 10'h3a0;
        mem[344] = 10'h32e;
        mem[345] = 10'h2a8;
        mem[346] = 10'h1ca;
        mem[347] = 10'h194;
        mem[348] = 10'h2b8;
        mem[349] = 10'h0dd;
        mem[350] = 10'h3f1;
        mem[351] = 10'h031;
        mem[352] = 10'h39d;
        mem[353] = 10'h026;
        mem[354] = 10'h244;
        mem[355] = 10'h02d;
        mem[356] = 10'h117;
        mem[357] = 10'h370;
        mem[358] = 10'h22d;
        mem[359] = 10'h2ea;
        mem[360] = 10'h165;
        mem[361] = 10'h115;
        mem[362] = 10'h167;
        mem[363] = 10'h3f4;
        mem[364] = 10'h0df;
        mem[365] = 10'h34f;
        mem[366] = 10'h380;
        mem[367] = 10'h1c3;
        mem[368] = 10'h0c8;
        mem[369] = 10'h3eb;
        mem[370] = 10'h325;
        mem[371] = 10'h051;
        mem[372] = 10'h1d2;
        mem[373] = 10'h13b;
        mem[374] = 10'h308;
        mem[375] = 10'h2ce;
        mem[376] = 10'h2b4;
        mem[377] = 10'h274;
        mem[378] = 10'h0a6;
        mem[379] = 10'h3e7;
        mem[380] = 10'h200;
        mem[381] = 10'h219;
        mem[382] = 10'h096;
        mem[383] = 10'h30f;
        mem[384] = 10'h177;
        mem[385] = 10'h09c;
        mem[386] = 10'h236;
        mem[387] = 10'h069;
        mem[388] = 10'h0d0;
        mem[389] = 10'h281;
        mem[390] = 10'h2e7;
        mem[391] = 10'h3b8;
        mem[392] = 10'h19a;
        mem[393] = 10'h235;
        mem[394] = 10'h122;
        mem[395] = 10'h20d;
        mem[396] = 10'h37b;
        mem[397] = 10'h091;
        mem[398] = 10'h3ba;
        mem[399] = 10'h362;
        mem[400] = 10'h2be;
        mem[401] = 10'h1b9;
        mem[402] = 10'h1f1;
        mem[403] = 10'h03d;
        mem[404] = 10'h29d;
        mem[405] = 10'h23a;
        mem[406] = 10'h296;
        mem[407] = 10'h21a;
        mem[408] = 10'h149;
        mem[409] = 10'h3ee;
        mem[410] = 10'h088;
        mem[411] = 10'h3e0;
        mem[412] = 10'h365;
        mem[413] = 10'h1cc;
        mem[414] = 10'h10d;
        mem[415] = 10'h1df;
        mem[416] = 10'h063;
        mem[417] = 10'h253;
        mem[418] = 10'h320;
        mem[419] = 10'h31e;
        mem[420] = 10'h2f3;
        mem[421] = 10'h08a;
        mem[422] = 10'h3d4;
        mem[423] = 10'h345;
        mem[424] = 10'h04c;
        mem[425] = 10'h09d;
        mem[426] = 10'h263;
        mem[427] = 10'h397;
        mem[428] = 10'h3e8;
        mem[429] = 10'h0e8;
        mem[430] = 10'h1e4;
        mem[431] = 10'h15d;
        mem[432] = 10'h3db;
        mem[433] = 10'h040;
        mem[434] = 10'h35f;
        mem[435] = 10'h3b0;
        mem[436] = 10'h070;
        mem[437] = 10'h21c;
        mem[438] = 10'h04e;
        mem[439] = 10'h1ac;
        mem[440] = 10'h28c;
        mem[441] = 10'h2b6;
        mem[442] = 10'h19e;
        mem[443] = 10'h0ec;
        mem[444] = 10'h2f7;
        mem[445] = 10'h113;
        mem[446] = 10'h0c9;
        mem[447] = 10'h1ad;
        mem[448] = 10'h02f;
        mem[449] = 10'h37a;
        mem[450] = 10'h36f;
        mem[451] = 10'h2dc;
        mem[452] = 10'h2eb;
        mem[453] = 10'h180;
        mem[454] = 10'h042;
        mem[455] = 10'h284;
        mem[456] = 10'h38d;
        mem[457] = 10'h25f;
        mem[458] = 10'h05d;
        mem[459] = 10'h1a9;
        mem[460] = 10'h257;
        mem[461] = 10'h2e3;
        mem[462] = 10'h24d;
        mem[463] = 10'h372;
        mem[464] = 10'h1e9;
        mem[465] = 10'h3d0;
        mem[466] = 10'h030;
        mem[467] = 10'h332;
        mem[468] = 10'h0c2;
        mem[469] = 10'h3cc;
        mem[470] = 10'h085;
        mem[471] = 10'h2c5;
        mem[472] = 10'h1ae;
        mem[473] = 10'h2a5;
        mem[474] = 10'h06f;
        mem[475] = 10'h2fd;
        mem[476] = 10'h2ae;
        mem[477] = 10'h2fb;
        mem[478] = 10'h256;
        mem[479] = 10'h282;
        mem[480] = 10'h373;
        mem[481] = 10'h1f8;
        mem[482] = 10'h379;
        mem[483] = 10'h17c;
        mem[484] = 10'h0f6;
        mem[485] = 10'h3bc;
        mem[486] = 10'h13e;
        mem[487] = 10'h3b7;
        mem[488] = 10'h271;
        mem[489] = 10'h3cf;
        mem[490] = 10'h19c;
        mem[491] = 10'h13c;
        mem[492] = 10'h25b;
        mem[493] = 10'h10e;
        mem[494] = 10'h0cc;
        mem[495] = 10'h1e1;
        mem[496] = 10'h0cb;
        mem[497] = 10'h2c4;
        mem[498] = 10'h377;
        mem[499] = 10'h38e;
        mem[500] = 10'h074;
        mem[501] = 10'h2a7;
        mem[502] = 10'h1c7;
        mem[503] = 10'h1f7;
        mem[504] = 10'h240;
        mem[505] = 10'h28b;
        mem[506] = 10'h1db;
        mem[507] = 10'h353;
        mem[508] = 10'h08f;
        mem[509] = 10'h29a;
        mem[510] = 10'h2c7;
        mem[511] = 10'h15c;
        mem[512] = 10'h3e3;
        mem[513] = 10'h1d9;
        mem[514] = 10'h1d5;
        mem[515] = 10'h2ac;
        mem[516] = 10'h22a;
        mem[517] = 10'h243;
        mem[518] = 10'h16e;
        mem[519] = 10'h214;
        mem[520] = 10'h0b8;
        mem[521] = 10'h36a;
        mem[522] = 10'h391;
        mem[523] = 10'h033;
        mem[524] = 10'h123;
        mem[525] = 10'h374;
        mem[526] = 10'h1e0;
        mem[527] = 10'h307;
        mem[528] = 10'h258;
        mem[529] = 10'h22b;
        mem[530] = 10'h216;
        mem[531] = 10'h2a6;
        mem[532] = 10'h0e1;
        mem[533] = 10'h196;
        mem[534] = 10'h0e4;
        mem[535] = 10'h3ff;
        mem[536] = 10'h2c6;
        mem[537] = 10'h0ba;
        mem[538] = 10'h3a2;
        mem[539] = 10'h38c;
        mem[540] = 10'h161;
        mem[541] = 10'h358;
        mem[542] = 10'h00e;
        mem[543] = 10'h06b;
        mem[544] = 10'h1cb;
        mem[545] = 10'h31c;
        mem[546] = 10'h3ca;
        mem[547] = 10'h023;
        mem[548] = 10'h3c3;
        mem[549] = 10'h24b;
        mem[550] = 10'h1c4;
        mem[551] = 10'h0eb;
        mem[552] = 10'h028;
        mem[553] = 10'h29c;
        mem[554] = 10'h0ab;
        mem[555] = 10'h1ef;
        mem[556] = 10'h0d4;
        mem[557] = 10'h049;
        mem[558] = 10'h2d5;
        mem[559] = 10'h139;
        mem[560] = 10'h22c;
        mem[561] = 10'h392;
        mem[562] = 10'h152;
        mem[563] = 10'h1ea;
        mem[564] = 10'h302;
        mem[565] = 10'h209;
        mem[566] = 10'h262;
        mem[567] = 10'h3f3;
        mem[568] = 10'h2f4;
        mem[569] = 10'h27d;
        mem[570] = 10'h335;
        mem[571] = 10'h2f1;
        mem[572] = 10'h130;
        mem[573] = 10'h338;
        mem[574] = 10'h0f9;
        mem[575] = 10'h2a3;
        mem[576] = 10'h12a;
        mem[577] = 10'h2a4;
        mem[578] = 10'h073;
        mem[579] = 10'h111;
        mem[580] = 10'h3a7;
        mem[581] = 10'h386;
        mem[582] = 10'h2e4;
        mem[583] = 10'h2f6;
        mem[584] = 10'h1c9;
        mem[585] = 10'h38a;
        mem[586] = 10'h2d8;
        mem[587] = 10'h341;
        mem[588] = 10'h0b6;
        mem[589] = 10'h05a;
        mem[590] = 10'h17f;
        mem[591] = 10'h037;
        mem[592] = 10'h29f;
        mem[593] = 10'h2fa;
        mem[594] = 10'h03b;
        mem[595] = 10'h00f;
        mem[596] = 10'h238;
        mem[597] = 10'h37f;
        mem[598] = 10'h265;
        mem[599] = 10'h169;
        mem[600] = 10'h09b;
        mem[601] = 10'h3c8;
        mem[602] = 10'h163;
        mem[603] = 10'h3fa;
        mem[604] = 10'h385;
        mem[605] = 10'h1b7;
        mem[606] = 10'h0f0;
        mem[607] = 10'h30d;
        mem[608] = 10'h035;
        mem[609] = 10'h067;
        mem[610] = 10'h1eb;
        mem[611] = 10'h280;
        mem[612] = 10'h3a9;
        mem[613] = 10'h245;
        mem[614] = 10'h0e5;
        mem[615] = 10'h311;
        mem[616] = 10'h141;
        mem[617] = 10'h22e;
        mem[618] = 10'h24c;
        mem[619] = 10'h247;
        mem[620] = 10'h28d;
        mem[621] = 10'h097;
        mem[622] = 10'h293;
        mem[623] = 10'h3c5;
        mem[624] = 10'h135;
        mem[625] = 10'h2fc;
        mem[626] = 10'h378;
        mem[627] = 10'h16d;
        mem[628] = 10'h1cf;
        mem[629] = 10'h198;
        mem[630] = 10'h317;
        mem[631] = 10'h05e;
        mem[632] = 10'h0ca;
        mem[633] = 10'h2ca;
        mem[634] = 10'h212;
        mem[635] = 10'h075;
        mem[636] = 10'h3c9;
        mem[637] = 10'h17d;
        mem[638] = 10'h26c;
        mem[639] = 10'h07f;
        mem[640] = 10'h269;
        mem[641] = 10'h2db;
        mem[642] = 10'h1aa;
        mem[643] = 10'h25c;
        mem[644] = 10'h190;
        mem[645] = 10'h3f7;
        mem[646] = 10'h292;
        mem[647] = 10'h129;
        mem[648] = 10'h1da;
        mem[649] = 10'h30b;
        mem[650] = 10'h26e;
        mem[651] = 10'h384;
        mem[652] = 10'h090;
        mem[653] = 10'h105;
        mem[654] = 10'h0be;
        mem[655] = 10'h254;
        mem[656] = 10'h188;
        mem[657] = 10'h259;
        mem[658] = 10'h19f;
        mem[659] = 10'h018;
        mem[660] = 10'h012;
        mem[661] = 10'h3cb;
        mem[662] = 10'h2ef;
        mem[663] = 10'h39b;
        mem[664] = 10'h0d5;
        mem[665] = 10'h2f0;
        mem[666] = 10'h354;
        mem[667] = 10'h28a;
        mem[668] = 10'h2b2;
        mem[669] = 10'h0b1;
        mem[670] = 10'h343;
        mem[671] = 10'h1e3;
        mem[672] = 10'h221;
        mem[673] = 10'h1b4;
        mem[674] = 10'h100;
        mem[675] = 10'h089;
        mem[676] = 10'h12b;
        mem[677] = 10'h20b;
        mem[678] = 10'h3e6;
        mem[679] = 10'h23f;
        mem[680] = 10'h275;
        mem[681] = 10'h35a;
        mem[682] = 10'h083;
        mem[683] = 10'h1bd;
        mem[684] = 10'h315;
        mem[685] = 10'h37c;
        mem[686] = 10'h12f;
        mem[687] = 10'h10a;
        mem[688] = 10'h052;
        mem[689] = 10'h208;
        mem[690] = 10'h0dc;
        mem[691] = 10'h095;
        mem[692] = 10'h002;
        mem[693] = 10'h04d;
        mem[694] = 10'h025;
        mem[695] = 10'h153;
        mem[696] = 10'h0cf;
        mem[697] = 10'h175;
        mem[698] = 10'h077;
        mem[699] = 10'h34b;
        mem[700] = 10'h14c;
        mem[701] = 10'h101;
        mem[702] = 10'h0a1;
        mem[703] = 10'h0d9;
        mem[704] = 10'h30c;
        mem[705] = 10'h3fd;
        mem[706] = 10'h0fb;
        mem[707] = 10'h3f9;
        mem[708] = 10'h106;
        mem[709] = 10'h387;
        mem[710] = 10'h12c;
        mem[711] = 10'h0ee;
        mem[712] = 10'h0db;
        mem[713] = 10'h1e8;
        mem[714] = 10'h2e8;
        mem[715] = 10'h3f2;
        mem[716] = 10'h2d3;
        mem[717] = 10'h3ce;
        mem[718] = 10'h30a;
        mem[719] = 10'h0b0;
        mem[720] = 10'h03e;
        mem[721] = 10'h1c0;
        mem[722] = 10'h398;
        mem[723] = 10'h327;
        mem[724] = 10'h283;
        mem[725] = 10'h034;
        mem[726] = 10'h1be;
        mem[727] = 10'h019;
        mem[728] = 10'h185;
        mem[729] = 10'h355;
        mem[730] = 10'h134;
        mem[731] = 10'h036;
        mem[732] = 10'h202;
        mem[733] = 10'h2d9;
        mem[734] = 10'h01b;
        mem[735] = 10'h102;
        mem[736] = 10'h06e;
        mem[737] = 10'h38b;
        mem[738] = 10'h191;
        mem[739] = 10'h076;
        mem[740] = 10'h399;
        mem[741] = 10'h126;
        mem[742] = 10'h1bc;
        mem[743] = 10'h043;
        mem[744] = 10'h156;
        mem[745] = 10'h087;
        mem[746] = 10'h160;
        mem[747] = 10'h0c5;
        mem[748] = 10'h022;
        mem[749] = 10'h1bf;
        mem[750] = 10'h26a;
        mem[751] = 10'h0de;
        mem[752] = 10'h33b;
        mem[753] = 10'h326;
        mem[754] = 10'h2c8;
        mem[755] = 10'h0a7;
        mem[756] = 10'h066;
        mem[757] = 10'h2fe;
        mem[758] = 10'h0b2;
        mem[759] = 10'h02a;
        mem[760] = 10'h2dd;
        mem[761] = 10'h1d3;
        mem[762] = 10'h3da;
        mem[763] = 10'h36c;
        mem[764] = 10'h04b;
        mem[765] = 10'h011;
        mem[766] = 10'h1ee;
        mem[767] = 10'h0ef;
        mem[768] = 10'h1ce;
        mem[769] = 10'h17b;
        mem[770] = 10'h1fa;
        mem[771] = 10'h295;
        mem[772] = 10'h0bf;
        mem[773] = 10'h12e;
        mem[774] = 10'h14d;
        mem[775] = 10'h31d;
        mem[776] = 10'h2df;
        mem[777] = 10'h0d7;
        mem[778] = 10'h055;
        mem[779] = 10'h394;
        mem[780] = 10'h1d1;
        mem[781] = 10'h289;
        mem[782] = 10'h01e;
        mem[783] = 10'h321;
        mem[784] = 10'h147;
        mem[785] = 10'h14a;
        mem[786] = 10'h047;
        mem[787] = 10'h34a;
        mem[788] = 10'h32b;
        mem[789] = 10'h3e2;
        mem[790] = 10'h21b;
        mem[791] = 10'h1e5;
        mem[792] = 10'h0aa;
        mem[793] = 10'h310;
        mem[794] = 10'h261;
        mem[795] = 10'h1c5;
        mem[796] = 10'h299;
        mem[797] = 10'h107;
        mem[798] = 10'h346;
        mem[799] = 10'h0e7;
        mem[800] = 10'h39c;
        mem[801] = 10'h2ab;
        mem[802] = 10'h2b7;
        mem[803] = 10'h3bf;
        mem[804] = 10'h13f;
        mem[805] = 10'h395;
        mem[806] = 10'h312;
        mem[807] = 10'h15b;
        mem[808] = 10'h1cd;
        mem[809] = 10'h2d1;
        mem[810] = 10'h148;
        mem[811] = 10'h229;
        mem[812] = 10'h3e4;
        mem[813] = 10'h290;
        mem[814] = 10'h0f8;
        mem[815] = 10'h1bb;
        mem[816] = 10'h068;
        mem[817] = 10'h1ec;
        mem[818] = 10'h13a;
        mem[819] = 10'h1fd;
        mem[820] = 10'h1dd;
        mem[821] = 10'h195;
        mem[822] = 10'h1e7;
        mem[823] = 10'h104;
        mem[824] = 10'h23e;
        mem[825] = 10'h137;
        mem[826] = 10'h121;
        mem[827] = 10'h1b1;
        mem[828] = 10'h1d7;
        mem[829] = 10'h0fa;
        mem[830] = 10'h3d7;
        mem[831] = 10'h288;
        mem[832] = 10'h2af;
        mem[833] = 10'h3b5;
        mem[834] = 10'h199;
        mem[835] = 10'h182;
        mem[836] = 10'h27a;
        mem[837] = 10'h3d2;
        mem[838] = 10'h18b;
        mem[839] = 10'h09e;
        mem[840] = 10'h3aa;
        mem[841] = 10'h1dc;
        mem[842] = 10'h20a;
        mem[843] = 10'h1d0;
        mem[844] = 10'h092;
        mem[845] = 10'h2c0;
        mem[846] = 10'h222;
        mem[847] = 10'h36b;
        mem[848] = 10'h1f3;
        mem[849] = 10'h127;
        mem[850] = 10'h0d1;
        mem[851] = 10'h252;
        mem[852] = 10'h16a;
        mem[853] = 10'h00c;
        mem[854] = 10'h27f;
        mem[855] = 10'h05c;
        mem[856] = 10'h2e6;
        mem[857] = 10'h30e;
        mem[858] = 10'h2a9;
        mem[859] = 10'h02c;
        mem[860] = 10'h082;
        mem[861] = 10'h364;
        mem[862] = 10'h05f;
        mem[863] = 10'h04a;
        mem[864] = 10'h3c1;
        mem[865] = 10'h116;
        mem[866] = 10'h2f8;
        mem[867] = 10'h3e9;
        mem[868] = 10'h231;
        mem[869] = 10'h15f;
        mem[870] = 10'h3a3;
        mem[871] = 10'h211;
        mem[872] = 10'h31b;
        mem[873] = 10'h388;
        mem[874] = 10'h064;
        mem[875] = 10'h304;
        mem[876] = 10'h23b;
        mem[877] = 10'h3ed;
        mem[878] = 10'h322;
        mem[879] = 10'h041;
        mem[880] = 10'h309;
        mem[881] = 10'h35b;
        mem[882] = 10'h3ae;
        mem[883] = 10'h09f;
        mem[884] = 10'h3ec;
        mem[885] = 10'h166;
        mem[886] = 10'h1f6;
        mem[887] = 10'h330;
        mem[888] = 10'h0d8;
        mem[889] = 10'h32c;
        mem[890] = 10'h32d;
        mem[891] = 10'h0fc;
        mem[892] = 10'h21d;
        mem[893] = 10'h29b;
        mem[894] = 10'h218;
        mem[895] = 10'h2ec;
        mem[896] = 10'h010;
        mem[897] = 10'h197;
        mem[898] = 10'h2cb;
        mem[899] = 10'h279;
        mem[900] = 10'h203;
        mem[901] = 10'h005;
        mem[902] = 10'h08c;
        mem[903] = 10'h3fe;
        mem[904] = 10'h14f;
        mem[905] = 10'h0bd;
        mem[906] = 10'h3b9;
        mem[907] = 10'h11a;
        mem[908] = 10'h164;
        mem[909] = 10'h120;
        mem[910] = 10'h227;
        mem[911] = 10'h3fb;
        mem[912] = 10'h3ef;
        mem[913] = 10'h0f2;
        mem[914] = 10'h242;
        mem[915] = 10'h0b3;
        mem[916] = 10'h340;
        mem[917] = 10'h3c0;
        mem[918] = 10'h33d;
        mem[919] = 10'h382;
        mem[920] = 10'h224;
        mem[921] = 10'h3ea;
        mem[922] = 10'h059;
        mem[923] = 10'h029;
        mem[924] = 10'h004;
        mem[925] = 10'h225;
        mem[926] = 10'h0e9;
        mem[927] = 10'h07b;
        mem[928] = 10'h349;
        mem[929] = 10'h133;
        mem[930] = 10'h03f;
        mem[931] = 10'h046;
        mem[932] = 10'h0fd;
        mem[933] = 10'h2e5;
        mem[934] = 10'h336;
        mem[935] = 10'h0c3;
        mem[936] = 10'h2e1;
        mem[937] = 10'h33f;
        mem[938] = 10'h25e;
        mem[939] = 10'h056;
        mem[940] = 10'h2d0;
        mem[941] = 10'h14e;
        mem[942] = 10'h03c;
        mem[943] = 10'h3b2;
        mem[944] = 10'h16f;
        mem[945] = 10'h178;
        mem[946] = 10'h3b6;
        mem[947] = 10'h1f9;
        mem[948] = 10'h3a8;
        mem[949] = 10'h0ea;
        mem[950] = 10'h1b5;
        mem[951] = 10'h154;
        mem[952] = 10'h35c;
        mem[953] = 10'h2b0;
        mem[954] = 10'h233;
        mem[955] = 10'h0ad;
        mem[956] = 10'h226;
        mem[957] = 10'h23d;
        mem[958] = 10'h2c2;
        mem[959] = 10'h2ff;
        mem[960] = 10'h050;
        mem[961] = 10'h291;
        mem[962] = 10'h32a;
        mem[963] = 10'h368;
        mem[964] = 10'h170;
        mem[965] = 10'h2bc;
        mem[966] = 10'h1b3;
        mem[967] = 10'h062;
        mem[968] = 10'h390;
        mem[969] = 10'h18c;
        mem[970] = 10'h204;
        mem[971] = 10'h151;
        mem[972] = 10'h109;
        mem[973] = 10'h01a;
        mem[974] = 10'h3d3;
        mem[975] = 10'h3dc;
        mem[976] = 10'h21f;
        mem[977] = 10'h0a2;
        mem[978] = 10'h3ad;
        mem[979] = 10'h04f;
        mem[980] = 10'h110;
        mem[981] = 10'h223;
        mem[982] = 10'h1e6;
        mem[983] = 10'h11d;
        mem[984] = 10'h1a5;
        mem[985] = 10'h18d;
        mem[986] = 10'h080;
        mem[987] = 10'h303;
        mem[988] = 10'h234;
        mem[989] = 10'h0ed;
        mem[990] = 10'h0c0;
        mem[991] = 10'h0bb;
        mem[992] = 10'h1a0;
        mem[993] = 10'h081;
        mem[994] = 10'h33c;
        mem[995] = 10'h0da;
        mem[996] = 10'h11f;
        mem[997] = 10'h344;
        mem[998] = 10'h2a1;
        mem[999] = 10'h39a;
        mem[1000] = 10'h2d2;
        mem[1001] = 10'h08b;
        mem[1002] = 10'h0bc;
        mem[1003] = 10'h03a;
        mem[1004] = 10'h2cd;
        mem[1005] = 10'h06c;
        mem[1006] = 10'h2b1;
        mem[1007] = 10'h270;
        mem[1008] = 10'h1c8;
        mem[1009] = 10'h015;
        mem[1010] = 10'h1f2;
        mem[1011] = 10'h0e3;
        mem[1012] = 10'h286;
        mem[1013] = 10'h0e2;
        mem[1014] = 10'h2b5;
        mem[1015] = 10'h181;
        mem[1016] = 10'h3bb;
        mem[1017] = 10'h2c3;
        mem[1018] = 10'h1fb;
        mem[1019] = 10'h331;
        mem[1020] = 10'h1a7;
        mem[1021] = 10'h24a;
        mem[1022] = 10'h287;
        mem[1023] = 10'h3df;
    end
endmodule

module odo_sbox_large3(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    (* ram_style = "block" *) reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h390;
        mem[1] = 10'h394;
        mem[2] = 10'h078;
        mem[3] = 10'h2da;
        mem[4] = 10'h2fc;
        mem[5] = 10'h205;
        mem[6] = 10'h29d;
        mem[7] = 10'h2a3;
        mem[8] = 10'h07a;
        mem[9] = 10'h1ef;
        mem[10] = 10'h286;
        mem[11] = 10'h195;
        mem[12] = 10'h109;
        mem[13] = 10'h083;
        mem[14] = 10'h005;
        mem[15] = 10'h38c;
        mem[16] = 10'h0a4;
        mem[17] = 10'h179;
        mem[18] = 10'h32a;
        mem[19] = 10'h142;
        mem[20] = 10'h379;
        mem[21] = 10'h3bb;
        mem[22] = 10'h14a;
        mem[23] = 10'h3bf;
        mem[24] = 10'h3bc;
        mem[25] = 10'h20e;
        mem[26] = 10'h336;
        mem[27] = 10'h13e;
        mem[28] = 10'h02a;
        mem[29] = 10'h17c;
        mem[30] = 10'h149;
        mem[31] = 10'h271;
        mem[32] = 10'h2cd;
        mem[33] = 10'h141;
        mem[34] = 10'h054;
        mem[35] = 10'h384;
        mem[36] = 10'h105;
        mem[37] = 10'h2df;
        mem[38] = 10'h395;
        mem[39] = 10'h244;
        mem[40] = 10'h03a;
        mem[41] = 10'h383;
        mem[42] = 10'h3d8;
        mem[43] = 10'h39d;
        mem[44] = 10'h114;
        mem[45] = 10'h345;
        mem[46] = 10'h131;
        mem[47] = 10'h280;
        mem[48] = 10'h3f1;
        mem[49] = 10'h1ba;
        mem[50] = 10'h00c;
        mem[51] = 10'h312;
        mem[52] = 10'h307;
        mem[53] = 10'h039;
        mem[54] = 10'h18f;
        mem[55] = 10'h05c;
        mem[56] = 10'h01d;
        mem[57] = 10'h09b;
        mem[58] = 10'h342;
        mem[59] = 10'h2d6;
        mem[60] = 10'h36f;
        mem[61] = 10'h3e4;
        mem[62] = 10'h3d0;
        mem[63] = 10'h143;
        mem[64] = 10'h377;
        mem[65] = 10'h253;
        mem[66] = 10'h0ab;
        mem[67] = 10'h100;
        mem[68] = 10'h364;
        mem[69] = 10'h10e;
        mem[70] = 10'h0b4;
        mem[71] = 10'h3f4;
        mem[72] = 10'h2a5;
        mem[73] = 10'h251;
        mem[74] = 10'h2d0;
        mem[75] = 10'h020;
        mem[76] = 10'h0ad;
        mem[77] = 10'h353;
        mem[78] = 10'h037;
        mem[79] = 10'h025;
        mem[80] = 10'h2ff;
        mem[81] = 10'h003;
        mem[82] = 10'h266;
        mem[83] = 10'h33b;
        mem[84] = 10'h137;
        mem[85] = 10'h2b1;
        mem[86] = 10'h265;
        mem[87] = 10'h11c;
        mem[88] = 10'h1a8;
        mem[89] = 10'h3bd;
        mem[90] = 10'h05d;
        mem[91] = 10'h106;
        mem[92] = 10'h208;
        mem[93] = 10'h375;
        mem[94] = 10'h086;
        mem[95] = 10'h3e0;
        mem[96] = 10'h2ea;
        mem[97] = 10'h181;
        mem[98] = 10'h3a7;
        mem[99] = 10'h339;
        mem[100] = 10'h0a0;
        mem[101] = 10'h156;
        mem[102] = 10'h372;
        mem[103] = 10'h258;
        mem[104] = 10'h215;
        mem[105] = 10'h3de;
        mem[106] = 10'h1f1;
        mem[107] = 10'h295;
        mem[108] = 10'h28e;
        mem[109] = 10'h3c4;
        mem[110] = 10'h255;
        mem[111] = 10'h34c;
        mem[112] = 10'h1b3;
        mem[113] = 10'h190;
        mem[114] = 10'h016;
        mem[115] = 10'h0b3;
        mem[116] = 10'h05f;
        mem[117] = 10'h1ce;
        mem[118] = 10'h168;
        mem[119] = 10'h3c0;
        mem[120] = 10'h02f;
        mem[121] = 10'h187;
        mem[122] = 10'h2c9;
        mem[123] = 10'h148;
        mem[124] = 10'h310;
        mem[125] = 10'h3df;
        mem[126] = 10'h16e;
        mem[127] = 10'h32b;
        mem[128] = 10'h0a2;
        mem[129] = 10'h2f5;
        mem[130] = 10'h27a;
        mem[131] = 10'h033;
        mem[132] = 10'h0ac;
        mem[133] = 10'h22a;
        mem[134] = 10'h2ad;
        mem[135] = 10'h044;
        mem[136] = 10'h3eb;
        mem[137] = 10'h370;
        mem[138] = 10'h08c;
        mem[139] = 10'h14f;
        mem[140] = 10'h071;
        mem[141] = 10'h3a0;
        mem[142] = 10'h099;
        mem[143] = 10'h1c4;
        mem[144] = 10'h18a;
        mem[145] = 10'h1cb;
        mem[146] = 10'h2c4;
        mem[147] = 10'h2a2;
        mem[148] = 10'h3d7;
        mem[149] = 10'h104;
        mem[150] = 10'h002;
        mem[151] = 10'h038;
        mem[152] = 10'h206;
        mem[153] = 10'h3b1;
        mem[154] = 10'h3af;
        mem[155] = 10'h3e9;
        mem[156] = 10'h093;
        mem[157] = 10'h1ea;
        mem[158] = 10'h25b;
        mem[159] = 10'h13a;
        mem[160] = 10'h39c;
        mem[161] = 10'h33f;
        mem[162] = 10'h39a;
        mem[163] = 10'h3ce;
        mem[164] = 10'h37f;
        mem[165] = 10'h20b;
        mem[166] = 10'h2c5;
        mem[167] = 10'h347;
        mem[168] = 10'h045;
        mem[169] = 10'h33e;
        mem[170] = 10'h10d;
        mem[171] = 10'h3fa;
        mem[172] = 10'h37d;
        mem[173] = 10'h04a;
        mem[174] = 10'h21f;
        mem[175] = 10'h069;
        mem[176] = 10'h225;
        mem[177] = 10'h01f;
        mem[178] = 10'h00d;
        mem[179] = 10'h0b2;
        mem[180] = 10'h283;
        mem[181] = 10'h21d;
        mem[182] = 10'h09d;
        mem[183] = 10'h06d;
        mem[184] = 10'h2cb;
        mem[185] = 10'h20c;
        mem[186] = 10'h33c;
        mem[187] = 10'h1ed;
        mem[188] = 10'h018;
        mem[189] = 10'h174;
        mem[190] = 10'h027;
        mem[191] = 10'h1ab;
        mem[192] = 10'h298;
        mem[193] = 10'h0e2;
        mem[194] = 10'h065;
        mem[195] = 10'h360;
        mem[196] = 10'h09f;
        mem[197] = 10'h267;
        mem[198] = 10'h315;
        mem[199] = 10'h02b;
        mem[200] = 10'h2c6;
        mem[201] = 10'h162;
        mem[202] = 10'h119;
        mem[203] = 10'h222;
        mem[204] = 10'h1d2;
        mem[205] = 10'h367;
        mem[206] = 10'h0da;
        mem[207] = 10'h210;
        mem[208] = 10'h14b;
        mem[209] = 10'h3e8;
        mem[210] = 10'h31b;
        mem[211] = 10'h01e;
        mem[212] = 10'h277;
        mem[213] = 10'h1d6;
        mem[214] = 10'h2e5;
        mem[215] = 10'h10f;
        mem[216] = 10'h3aa;
        mem[217] = 10'h0c2;
        mem[218] = 10'h31f;
        mem[219] = 10'h311;
        mem[220] = 10'h1c7;
        mem[221] = 10'h24a;
        mem[222] = 10'h3d2;
        mem[223] = 10'h3f2;
        mem[224] = 10'h0ea;
        mem[225] = 10'h08f;
        mem[226] = 10'h1fd;
        mem[227] = 10'h1e0;
        mem[228] = 10'h3f6;
        mem[229] = 10'h055;
        mem[230] = 10'h2ee;
        mem[231] = 10'h392;
        mem[232] = 10'h031;
        mem[233] = 10'h0df;
        mem[234] = 10'h158;
        mem[235] = 10'h2ce;
        mem[236] = 10'h219;
        mem[237] = 10'h396;
        mem[238] = 10'h35a;
        mem[239] = 10'h128;
        mem[240] = 10'h1c0;
        mem[241] = 10'h0c9;
        mem[242] = 10'h028;
        mem[243] = 10'h332;
        mem[244] = 10'h2b0;
        mem[245] = 10'h19c;
        mem[246] = 10'h296;
        mem[247] = 10'h3b2;
        mem[248] = 10'h352;
        mem[249] = 10'h080;
        mem[250] = 10'h2f1;
        mem[251] = 10'h2a4;
        mem[252] = 10'h161;
        mem[253] = 10'h0ca;
        mem[254] = 10'h130;
        mem[255] = 10'h308;
        mem[256] = 10'h110;
        mem[257] = 10'h0ee;
        mem[258] = 10'h073;
        mem[259] = 10'h38a;
        mem[260] = 10'h01b;
        mem[261] = 10'h31d;
        mem[262] = 10'h035;
        mem[263] = 10'h124;
        mem[264] = 10'h261;
        mem[265] = 10'h1b5;
        mem[266] = 10'h282;
        mem[267] = 10'h05b;
        mem[268] = 10'h06f;
        mem[269] = 10'h28d;
        mem[270] = 10'h328;
        mem[271] = 10'h052;
        mem[272] = 10'h07f;
        mem[273] = 10'h0bd;
        mem[274] = 10'h2f7;
        mem[275] = 10'h3b0;
        mem[276] = 10'h0b1;
        mem[277] = 10'h20a;
        mem[278] = 10'h115;
        mem[279] = 10'h3ee;
        mem[280] = 10'h1da;
        mem[281] = 10'h1bc;
        mem[282] = 10'h2de;
        mem[283] = 10'h272;
        mem[284] = 10'h07e;
        mem[285] = 10'h0be;
        mem[286] = 10'h064;
        mem[287] = 10'h2a1;
        mem[288] = 10'h38f;
        mem[289] = 10'h0c7;
        mem[290] = 10'h1b1;
        mem[291] = 10'h111;
        mem[292] = 10'h082;
        mem[293] = 10'h11d;
        mem[294] = 10'h117;
        mem[295] = 10'h0fd;
        mem[296] = 10'h182;
        mem[297] = 10'h092;
        mem[298] = 10'h123;
        mem[299] = 10'h3fc;
        mem[300] = 10'h2e9;
        mem[301] = 10'h2f0;
        mem[302] = 10'h254;
        mem[303] = 10'h343;
        mem[304] = 10'h062;
        mem[305] = 10'h040;
        mem[306] = 10'h2d2;
        mem[307] = 10'h301;
        mem[308] = 10'h217;
        mem[309] = 10'h096;
        mem[310] = 10'h3c6;
        mem[311] = 10'h232;
        mem[312] = 10'h3cf;
        mem[313] = 10'h238;
        mem[314] = 10'h326;
        mem[315] = 10'h160;
        mem[316] = 10'h37b;
        mem[317] = 10'h306;
        mem[318] = 10'h197;
        mem[319] = 10'h368;
        mem[320] = 10'h2b2;
        mem[321] = 10'h391;
        mem[322] = 10'h0e6;
        mem[323] = 10'h39b;
        mem[324] = 10'h17f;
        mem[325] = 10'h170;
        mem[326] = 10'h27c;
        mem[327] = 10'h324;
        mem[328] = 10'h293;
        mem[329] = 10'h021;
        mem[330] = 10'h1f5;
        mem[331] = 10'h26f;
        mem[332] = 10'h2dd;
        mem[333] = 10'h2db;
        mem[334] = 10'h30a;
        mem[335] = 10'h3ed;
        mem[336] = 10'h15d;
        mem[337] = 10'h34b;
        mem[338] = 10'h0b5;
        mem[339] = 10'h366;
        mem[340] = 10'h010;
        mem[341] = 10'h14e;
        mem[342] = 10'h3f9;
        mem[343] = 10'h2d4;
        mem[344] = 10'h0ae;
        mem[345] = 10'h24b;
        mem[346] = 10'h369;
        mem[347] = 10'h3cc;
        mem[348] = 10'h0b6;
        mem[349] = 10'h1e1;
        mem[350] = 10'h0c4;
        mem[351] = 10'h37e;
        mem[352] = 10'h1d9;
        mem[353] = 10'h3ac;
        mem[354] = 10'h393;
        mem[355] = 10'h1d3;
        mem[356] = 10'h103;
        mem[357] = 10'h25a;
        mem[358] = 10'h14d;
        mem[359] = 10'h285;
        mem[360] = 10'h0cd;
        mem[361] = 10'h1f7;
        mem[362] = 10'h1ad;
        mem[363] = 10'h178;
        mem[364] = 10'h365;
        mem[365] = 10'h333;
        mem[366] = 10'h243;
        mem[367] = 10'h127;
        mem[368] = 10'h1c3;
        mem[369] = 10'h1b6;
        mem[370] = 10'h042;
        mem[371] = 10'h3f5;
        mem[372] = 10'h221;
        mem[373] = 10'h1e3;
        mem[374] = 10'h28c;
        mem[375] = 10'h07b;
        mem[376] = 10'h2a0;
        mem[377] = 10'h17e;
        mem[378] = 10'h3dc;
        mem[379] = 10'h157;
        mem[380] = 10'h218;
        mem[381] = 10'h338;
        mem[382] = 10'h0e4;
        mem[383] = 10'h357;
        mem[384] = 10'h36d;
        mem[385] = 10'h3e1;
        mem[386] = 10'h1e6;
        mem[387] = 10'h3b6;
        mem[388] = 10'h171;
        mem[389] = 10'h346;
        mem[390] = 10'h382;
        mem[391] = 10'h227;
        mem[392] = 10'h37c;
        mem[393] = 10'h28f;
        mem[394] = 10'h2d1;
        mem[395] = 10'h0e3;
        mem[396] = 10'h2cc;
        mem[397] = 10'h2dc;
        mem[398] = 10'h29c;
        mem[399] = 10'h146;
        mem[400] = 10'h165;
        mem[401] = 10'h04e;
        mem[402] = 10'h3f7;
        mem[403] = 10'h17d;
        mem[404] = 10'h11f;
        mem[405] = 10'h007;
        mem[406] = 10'h089;
        mem[407] = 10'h00b;
        mem[408] = 10'h18d;
        mem[409] = 10'h25d;
        mem[410] = 10'h303;
        mem[411] = 10'h2af;
        mem[412] = 10'h3ff;
        mem[413] = 10'h1eb;
        mem[414] = 10'h116;
        mem[415] = 10'h34f;
        mem[416] = 10'h389;
        mem[417] = 10'h085;
        mem[418] = 10'h013;
        mem[419] = 10'h380;
        mem[420] = 10'h2d3;
        mem[421] = 10'h0f2;
        mem[422] = 10'h3d3;
        mem[423] = 10'h1ac;
        mem[424] = 10'h06b;
        mem[425] = 10'h36b;
        mem[426] = 10'h223;
        mem[427] = 10'h1fe;
        mem[428] = 10'h0f4;
        mem[429] = 10'h314;
        mem[430] = 10'h214;
        mem[431] = 10'h1b4;
        mem[432] = 10'h3c2;
        mem[433] = 10'h166;
        mem[434] = 10'h133;
        mem[435] = 10'h2d5;
        mem[436] = 10'h3a4;
        mem[437] = 10'h19e;
        mem[438] = 10'h38e;
        mem[439] = 10'h04b;
        mem[440] = 10'h3ef;
        mem[441] = 10'h1a4;
        mem[442] = 10'h350;
        mem[443] = 10'h3f3;
        mem[444] = 10'h2bd;
        mem[445] = 10'h14c;
        mem[446] = 10'h0f0;
        mem[447] = 10'h049;
        mem[448] = 10'h2c7;
        mem[449] = 10'h061;
        mem[450] = 10'h1b8;
        mem[451] = 10'h234;
        mem[452] = 10'h1a0;
        mem[453] = 10'h26d;
        mem[454] = 10'h2e4;
        mem[455] = 10'h27e;
        mem[456] = 10'h1ff;
        mem[457] = 10'h358;
        mem[458] = 10'h356;
        mem[459] = 10'h361;
        mem[460] = 10'h0c0;
        mem[461] = 10'h1de;
        mem[462] = 10'h12c;
        mem[463] = 10'h011;
        mem[464] = 10'h03c;
        mem[465] = 10'h2c0;
        mem[466] = 10'h08a;
        mem[467] = 10'h23f;
        mem[468] = 10'h24c;
        mem[469] = 10'h1c1;
        mem[470] = 10'h32d;
        mem[471] = 10'h067;
        mem[472] = 10'h2ae;
        mem[473] = 10'h019;
        mem[474] = 10'h2bb;
        mem[475] = 10'h063;
        mem[476] = 10'h3a2;
        mem[477] = 10'h01a;
        mem[478] = 10'h275;
        mem[479] = 10'h2a7;
        mem[480] = 10'h017;
        mem[481] = 10'h297;
        mem[482] = 10'h23d;
        mem[483] = 10'h22f;
        mem[484] = 10'h348;
        mem[485] = 10'h077;
        mem[486] = 10'h0d1;
        mem[487] = 10'h136;
        mem[488] = 10'h3b4;
        mem[489] = 10'h3ea;
        mem[490] = 10'h102;
        mem[491] = 10'h33d;
        mem[492] = 10'h3a8;
        mem[493] = 10'h2c1;
        mem[494] = 10'h0cb;
        mem[495] = 10'h2ef;
        mem[496] = 10'h21c;
        mem[497] = 10'h2e2;
        mem[498] = 10'h0b8;
        mem[499] = 10'h385;
        mem[500] = 10'h1fc;
        mem[501] = 10'h129;
        mem[502] = 10'h320;
        mem[503] = 10'h126;
        mem[504] = 10'h186;
        mem[505] = 10'h006;
        mem[506] = 10'h1fa;
        mem[507] = 10'h3fb;
        mem[508] = 10'h145;
        mem[509] = 10'h0c6;
        mem[510] = 10'h1a3;
        mem[511] = 10'h281;
        mem[512] = 10'h163;
        mem[513] = 10'h292;
        mem[514] = 10'h1bd;
        mem[515] = 10'h29e;
        mem[516] = 10'h35d;
        mem[517] = 10'h21a;
        mem[518] = 10'h386;
        mem[519] = 10'h3ec;
        mem[520] = 10'h081;
        mem[521] = 10'h23c;
        mem[522] = 10'h0fa;
        mem[523] = 10'h262;
        mem[524] = 10'h08b;
        mem[525] = 10'h135;
        mem[526] = 10'h304;
        mem[527] = 10'h098;
        mem[528] = 10'h2fa;
        mem[529] = 10'h2b4;
        mem[530] = 10'h381;
        mem[531] = 10'h25f;
        mem[532] = 10'h07d;
        mem[533] = 10'h300;
        mem[534] = 10'h2f6;
        mem[535] = 10'h2c8;
        mem[536] = 10'h188;
        mem[537] = 10'h229;
        mem[538] = 10'h241;
        mem[539] = 10'h29b;
        mem[540] = 10'h23a;
        mem[541] = 10'h3d4;
        mem[542] = 10'h274;
        mem[543] = 10'h159;
        mem[544] = 10'h134;
        mem[545] = 10'h175;
        mem[546] = 10'h2c2;
        mem[547] = 10'h0d5;
        mem[548] = 10'h184;
        mem[549] = 10'h30b;
        mem[550] = 10'h0fe;
        mem[551] = 10'h3c8;
        mem[552] = 10'h235;
        mem[553] = 10'h25c;
        mem[554] = 10'h2bf;
        mem[555] = 10'h090;
        mem[556] = 10'h0e1;
        mem[557] = 10'h057;
        mem[558] = 10'h147;
        mem[559] = 10'h125;
        mem[560] = 10'h329;
        mem[561] = 10'h059;
        mem[562] = 10'h075;
        mem[563] = 10'h0aa;
        mem[564] = 10'h3db;
        mem[565] = 10'h249;
        mem[566] = 10'h08d;
        mem[567] = 10'h305;
        mem[568] = 10'h399;
        mem[569] = 10'h084;
        mem[570] = 10'h22c;
        mem[571] = 10'h2ca;
        mem[572] = 10'h25e;
        mem[573] = 10'h0bf;
        mem[574] = 10'h36c;
        mem[575] = 10'h0e5;
        mem[576] = 10'h0d3;
        mem[577] = 10'h30e;
        mem[578] = 10'h245;
        mem[579] = 10'h2e3;
        mem[580] = 10'h056;
        mem[581] = 10'h278;
        mem[582] = 10'h034;
        mem[583] = 10'h2be;
        mem[584] = 10'h199;
        mem[585] = 10'h3ca;
        mem[586] = 10'h28a;
        mem[587] = 10'h15f;
        mem[588] = 10'h378;
        mem[589] = 10'h371;
        mem[590] = 10'h1ae;
        mem[591] = 10'h070;
        mem[592] = 10'h202;
        mem[593] = 10'h0cc;
        mem[594] = 10'h1c9;
        mem[595] = 10'h0a5;
        mem[596] = 10'h1f4;
        mem[597] = 10'h3e6;
        mem[598] = 10'h2e6;
        mem[599] = 10'h26a;
        mem[600] = 10'h22d;
        mem[601] = 10'h240;
        mem[602] = 10'h06c;
        mem[603] = 10'h321;
        mem[604] = 10'h23e;
        mem[605] = 10'h327;
        mem[606] = 10'h30f;
        mem[607] = 10'h0f7;
        mem[608] = 10'h09e;
        mem[609] = 10'h2a8;
        mem[610] = 10'h1af;
        mem[611] = 10'h0f1;
        mem[612] = 10'h0ec;
        mem[613] = 10'h30c;
        mem[614] = 10'h176;
        mem[615] = 10'h374;
        mem[616] = 10'h1dc;
        mem[617] = 10'h1c8;
        mem[618] = 10'h001;
        mem[619] = 10'h1e4;
        mem[620] = 10'h39e;
        mem[621] = 10'h3fe;
        mem[622] = 10'h3ba;
        mem[623] = 10'h290;
        mem[624] = 10'h076;
        mem[625] = 10'h046;
        mem[626] = 10'h0b7;
        mem[627] = 10'h097;
        mem[628] = 10'h3b7;
        mem[629] = 10'h0fb;
        mem[630] = 10'h3d1;
        mem[631] = 10'h226;
        mem[632] = 10'h236;
        mem[633] = 10'h066;
        mem[634] = 10'h0ef;
        mem[635] = 10'h13d;
        mem[636] = 10'h16d;
        mem[637] = 10'h060;
        mem[638] = 10'h1dd;
        mem[639] = 10'h196;
        mem[640] = 10'h3b9;
        mem[641] = 10'h20f;
        mem[642] = 10'h164;
        mem[643] = 10'h3dd;
        mem[644] = 10'h172;
        mem[645] = 10'h207;
        mem[646] = 10'h38d;
        mem[647] = 10'h2e0;
        mem[648] = 10'h3cd;
        mem[649] = 10'h15a;
        mem[650] = 10'h318;
        mem[651] = 10'h014;
        mem[652] = 10'h23b;
        mem[653] = 10'h2a6;
        mem[654] = 10'h05a;
        mem[655] = 10'h2eb;
        mem[656] = 10'h27d;
        mem[657] = 10'h3b3;
        mem[658] = 10'h091;
        mem[659] = 10'h259;
        mem[660] = 10'h3a9;
        mem[661] = 10'h1f3;
        mem[662] = 10'h1df;
        mem[663] = 10'h2e7;
        mem[664] = 10'h0a7;
        mem[665] = 10'h012;
        mem[666] = 10'h0db;
        mem[667] = 10'h1f0;
        mem[668] = 10'h35b;
        mem[669] = 10'h3d6;
        mem[670] = 10'h287;
        mem[671] = 10'h36e;
        mem[672] = 10'h34d;
        mem[673] = 10'h322;
        mem[674] = 10'h387;
        mem[675] = 10'h24f;
        mem[676] = 10'h18b;
        mem[677] = 10'h309;
        mem[678] = 10'h26b;
        mem[679] = 10'h1e9;
        mem[680] = 10'h34e;
        mem[681] = 10'h1a5;
        mem[682] = 10'h39f;
        mem[683] = 10'h030;
        mem[684] = 10'h029;
        mem[685] = 10'h004;
        mem[686] = 10'h0a6;
        mem[687] = 10'h0a8;
        mem[688] = 10'h242;
        mem[689] = 10'h00a;
        mem[690] = 10'h04f;
        mem[691] = 10'h2e8;
        mem[692] = 10'h354;
        mem[693] = 10'h3cb;
        mem[694] = 10'h13f;
        mem[695] = 10'h230;
        mem[696] = 10'h1c2;
        mem[697] = 10'h113;
        mem[698] = 10'h0d4;
        mem[699] = 10'h2ec;
        mem[700] = 10'h237;
        mem[701] = 10'h29f;
        mem[702] = 10'h0d9;
        mem[703] = 10'h231;
        mem[704] = 10'h331;
        mem[705] = 10'h2b9;
        mem[706] = 10'h04c;
        mem[707] = 10'h11b;
        mem[708] = 10'h139;
        mem[709] = 10'h1ca;
        mem[710] = 10'h191;
        mem[711] = 10'h15e;
        mem[712] = 10'h2aa;
        mem[713] = 10'h3c3;
        mem[714] = 10'h3e3;
        mem[715] = 10'h1c6;
        mem[716] = 10'h000;
        mem[717] = 10'h1e2;
        mem[718] = 10'h0c3;
        mem[719] = 10'h35c;
        mem[720] = 10'h048;
        mem[721] = 10'h0a9;
        mem[722] = 10'h043;
        mem[723] = 10'h1ec;
        mem[724] = 10'h3a3;
        mem[725] = 10'h2f9;
        mem[726] = 10'h169;
        mem[727] = 10'h12e;
        mem[728] = 10'h3ad;
        mem[729] = 10'h183;
        mem[730] = 10'h36a;
        mem[731] = 10'h108;
        mem[732] = 10'h2e1;
        mem[733] = 10'h3fd;
        mem[734] = 10'h33a;
        mem[735] = 10'h27f;
        mem[736] = 10'h008;
        mem[737] = 10'h24d;
        mem[738] = 10'h047;
        mem[739] = 10'h2fb;
        mem[740] = 10'h3c7;
        mem[741] = 10'h1bb;
        mem[742] = 10'h140;
        mem[743] = 10'h2fd;
        mem[744] = 10'h05e;
        mem[745] = 10'h294;
        mem[746] = 10'h0fc;
        mem[747] = 10'h3e5;
        mem[748] = 10'h330;
        mem[749] = 10'h12a;
        mem[750] = 10'h1a6;
        mem[751] = 10'h0c1;
        mem[752] = 10'h20d;
        mem[753] = 10'h291;
        mem[754] = 10'h3ae;
        mem[755] = 10'h1f6;
        mem[756] = 10'h2c3;
        mem[757] = 10'h1cf;
        mem[758] = 10'h2b8;
        mem[759] = 10'h154;
        mem[760] = 10'h1f2;
        mem[761] = 10'h04d;
        mem[762] = 10'h1d4;
        mem[763] = 10'h323;
        mem[764] = 10'h3b8;
        mem[765] = 10'h239;
        mem[766] = 10'h0f8;
        mem[767] = 10'h248;
        mem[768] = 10'h03b;
        mem[769] = 10'h112;
        mem[770] = 10'h1aa;
        mem[771] = 10'h09c;
        mem[772] = 10'h12d;
        mem[773] = 10'h373;
        mem[774] = 10'h07c;
        mem[775] = 10'h32f;
        mem[776] = 10'h325;
        mem[777] = 10'h334;
        mem[778] = 10'h173;
        mem[779] = 10'h2b6;
        mem[780] = 10'h397;
        mem[781] = 10'h107;
        mem[782] = 10'h302;
        mem[783] = 10'h38b;
        mem[784] = 10'h31c;
        mem[785] = 10'h269;
        mem[786] = 10'h35e;
        mem[787] = 10'h198;
        mem[788] = 10'h153;
        mem[789] = 10'h273;
        mem[790] = 10'h247;
        mem[791] = 10'h0e0;
        mem[792] = 10'h0d8;
        mem[793] = 10'h316;
        mem[794] = 10'h058;
        mem[795] = 10'h138;
        mem[796] = 10'h212;
        mem[797] = 10'h120;
        mem[798] = 10'h10c;
        mem[799] = 10'h3da;
        mem[800] = 10'h01c;
        mem[801] = 10'h220;
        mem[802] = 10'h2b7;
        mem[803] = 10'h203;
        mem[804] = 10'h13c;
        mem[805] = 10'h22b;
        mem[806] = 10'h079;
        mem[807] = 10'h344;
        mem[808] = 10'h0af;
        mem[809] = 10'h1b2;
        mem[810] = 10'h0eb;
        mem[811] = 10'h0ed;
        mem[812] = 10'h16b;
        mem[813] = 10'h2ab;
        mem[814] = 10'h02e;
        mem[815] = 10'h1d7;
        mem[816] = 10'h276;
        mem[817] = 10'h194;
        mem[818] = 10'h3c5;
        mem[819] = 10'h122;
        mem[820] = 10'h12f;
        mem[821] = 10'h050;
        mem[822] = 10'h260;
        mem[823] = 10'h211;
        mem[824] = 10'h185;
        mem[825] = 10'h313;
        mem[826] = 10'h3e7;
        mem[827] = 10'h08e;
        mem[828] = 10'h233;
        mem[829] = 10'h053;
        mem[830] = 10'h0c5;
        mem[831] = 10'h023;
        mem[832] = 10'h264;
        mem[833] = 10'h27b;
        mem[834] = 10'h270;
        mem[835] = 10'h17a;
        mem[836] = 10'h3d5;
        mem[837] = 10'h0de;
        mem[838] = 10'h24e;
        mem[839] = 10'h1f9;
        mem[840] = 10'h2f3;
        mem[841] = 10'h009;
        mem[842] = 10'h341;
        mem[843] = 10'h101;
        mem[844] = 10'h121;
        mem[845] = 10'h2fe;
        mem[846] = 10'h03f;
        mem[847] = 10'h349;
        mem[848] = 10'h3a1;
        mem[849] = 10'h22e;
        mem[850] = 10'h151;
        mem[851] = 10'h3d9;
        mem[852] = 10'h06e;
        mem[853] = 10'h1ee;
        mem[854] = 10'h228;
        mem[855] = 10'h201;
        mem[856] = 10'h152;
        mem[857] = 10'h28b;
        mem[858] = 10'h094;
        mem[859] = 10'h21e;
        mem[860] = 10'h21b;
        mem[861] = 10'h3b5;
        mem[862] = 10'h0a1;
        mem[863] = 10'h17b;
        mem[864] = 10'h1a1;
        mem[865] = 10'h376;
        mem[866] = 10'h1fb;
        mem[867] = 10'h16c;
        mem[868] = 10'h095;
        mem[869] = 10'h167;
        mem[870] = 10'h0c8;
        mem[871] = 10'h088;
        mem[872] = 10'h024;
        mem[873] = 10'h2d8;
        mem[874] = 10'h3c1;
        mem[875] = 10'h02d;
        mem[876] = 10'h11a;
        mem[877] = 10'h279;
        mem[878] = 10'h16a;
        mem[879] = 10'h31a;
        mem[880] = 10'h30d;
        mem[881] = 10'h1cd;
        mem[882] = 10'h319;
        mem[883] = 10'h0f9;
        mem[884] = 10'h1b0;
        mem[885] = 10'h0d2;
        mem[886] = 10'h026;
        mem[887] = 10'h09a;
        mem[888] = 10'h1e8;
        mem[889] = 10'h26e;
        mem[890] = 10'h0f5;
        mem[891] = 10'h02c;
        mem[892] = 10'h00f;
        mem[893] = 10'h2f8;
        mem[894] = 10'h144;
        mem[895] = 10'h317;
        mem[896] = 10'h015;
        mem[897] = 10'h18c;
        mem[898] = 10'h388;
        mem[899] = 10'h0f3;
        mem[900] = 10'h3f8;
        mem[901] = 10'h0bc;
        mem[902] = 10'h37a;
        mem[903] = 10'h362;
        mem[904] = 10'h1e7;
        mem[905] = 10'h10b;
        mem[906] = 10'h26c;
        mem[907] = 10'h1a2;
        mem[908] = 10'h1d0;
        mem[909] = 10'h118;
        mem[910] = 10'h3ab;
        mem[911] = 10'h1c5;
        mem[912] = 10'h13b;
        mem[913] = 10'h263;
        mem[914] = 10'h351;
        mem[915] = 10'h0b0;
        mem[916] = 10'h2cf;
        mem[917] = 10'h022;
        mem[918] = 10'h355;
        mem[919] = 10'h1d5;
        mem[920] = 10'h16f;
        mem[921] = 10'h1d8;
        mem[922] = 10'h051;
        mem[923] = 10'h0e8;
        mem[924] = 10'h1a9;
        mem[925] = 10'h289;
        mem[926] = 10'h15b;
        mem[927] = 10'h2bc;
        mem[928] = 10'h132;
        mem[929] = 10'h0f6;
        mem[930] = 10'h3f0;
        mem[931] = 10'h1bf;
        mem[932] = 10'h041;
        mem[933] = 10'h0d7;
        mem[934] = 10'h1f8;
        mem[935] = 10'h224;
        mem[936] = 10'h31e;
        mem[937] = 10'h2f2;
        mem[938] = 10'h3a5;
        mem[939] = 10'h34a;
        mem[940] = 10'h3be;
        mem[941] = 10'h0e9;
        mem[942] = 10'h299;
        mem[943] = 10'h06a;
        mem[944] = 10'h150;
        mem[945] = 10'h1d1;
        mem[946] = 10'h200;
        mem[947] = 10'h19f;
        mem[948] = 10'h0dd;
        mem[949] = 10'h288;
        mem[950] = 10'h0d6;
        mem[951] = 10'h3c9;
        mem[952] = 10'h1e5;
        mem[953] = 10'h257;
        mem[954] = 10'h2ed;
        mem[955] = 10'h155;
        mem[956] = 10'h0ff;
        mem[957] = 10'h363;
        mem[958] = 10'h177;
        mem[959] = 10'h03e;
        mem[960] = 10'h209;
        mem[961] = 10'h250;
        mem[962] = 10'h1cc;
        mem[963] = 10'h19a;
        mem[964] = 10'h0d0;
        mem[965] = 10'h074;
        mem[966] = 10'h256;
        mem[967] = 10'h03d;
        mem[968] = 10'h11e;
        mem[969] = 10'h337;
        mem[970] = 10'h335;
        mem[971] = 10'h32e;
        mem[972] = 10'h10a;
        mem[973] = 10'h0ce;
        mem[974] = 10'h072;
        mem[975] = 10'h00e;
        mem[976] = 10'h2ac;
        mem[977] = 10'h0e7;
        mem[978] = 10'h036;
        mem[979] = 10'h068;
        mem[980] = 10'h0a3;
        mem[981] = 10'h35f;
        mem[982] = 10'h0bb;
        mem[983] = 10'h268;
        mem[984] = 10'h15c;
        mem[985] = 10'h1a7;
        mem[986] = 10'h032;
        mem[987] = 10'h2b3;
        mem[988] = 10'h3a6;
        mem[989] = 10'h359;
        mem[990] = 10'h1db;
        mem[991] = 10'h19b;
        mem[992] = 10'h180;
        mem[993] = 10'h284;
        mem[994] = 10'h213;
        mem[995] = 10'h19d;
        mem[996] = 10'h087;
        mem[997] = 10'h1b9;
        mem[998] = 10'h340;
        mem[999] = 10'h398;
        mem[1000] = 10'h2a9;
        mem[1001] = 10'h192;
        mem[1002] = 10'h252;
        mem[1003] = 10'h2d9;
        mem[1004] = 10'h1b7;
        mem[1005] = 10'h193;
        mem[1006] = 10'h3e2;
        mem[1007] = 10'h1be;
        mem[1008] = 10'h32c;
        mem[1009] = 10'h29a;
        mem[1010] = 10'h0b9;
        mem[1011] = 10'h204;
        mem[1012] = 10'h246;
        mem[1013] = 10'h0dc;
        mem[1014] = 10'h2d7;
        mem[1015] = 10'h2ba;
        mem[1016] = 10'h216;
        mem[1017] = 10'h2b5;
        mem[1018] = 10'h2f4;
        mem[1019] = 10'h12b;
        mem[1020] = 10'h189;
        mem[1021] = 10'h0cf;
        mem[1022] = 10'h0ba;
        mem[1023] = 10'h18e;
    end
endmodule

module odo_sbox_large4(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    (* ram_style = "block" *) reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h113;
        mem[1] = 10'h1a3;
        mem[2] = 10'h0f9;
        mem[3] = 10'h250;
        mem[4] = 10'h02f;
        mem[5] = 10'h1ca;
        mem[6] = 10'h0ba;
        mem[7] = 10'h363;
        mem[8] = 10'h037;
        mem[9] = 10'h0db;
        mem[10] = 10'h126;
        mem[11] = 10'h3ab;
        mem[12] = 10'h097;
        mem[13] = 10'h266;
        mem[14] = 10'h237;
        mem[15] = 10'h197;
        mem[16] = 10'h1a7;
        mem[17] = 10'h23d;
        mem[18] = 10'h2eb;
        mem[19] = 10'h371;
        mem[20] = 10'h367;
        mem[21] = 10'h252;
        mem[22] = 10'h1f3;
        mem[23] = 10'h0fa;
        mem[24] = 10'h2a9;
        mem[25] = 10'h392;
        mem[26] = 10'h077;
        mem[27] = 10'h3c2;
        mem[28] = 10'h2c5;
        mem[29] = 10'h272;
        mem[30] = 10'h1b3;
        mem[31] = 10'h036;
        mem[32] = 10'h07b;
        mem[33] = 10'h1e8;
        mem[34] = 10'h370;
        mem[35] = 10'h19f;
        mem[36] = 10'h2ff;
        mem[37] = 10'h3c0;
        mem[38] = 10'h1ec;
        mem[39] = 10'h222;
        mem[40] = 10'h3bb;
        mem[41] = 10'h093;
        mem[42] = 10'h0e8;
        mem[43] = 10'h046;
        mem[44] = 10'h29a;
        mem[45] = 10'h11f;
        mem[46] = 10'h25d;
        mem[47] = 10'h31e;
        mem[48] = 10'h368;
        mem[49] = 10'h191;
        mem[50] = 10'h092;
        mem[51] = 10'h1d1;
        mem[52] = 10'h1b4;
        mem[53] = 10'h159;
        mem[54] = 10'h234;
        mem[55] = 10'h090;
        mem[56] = 10'h2b9;
        mem[57] = 10'h175;
        mem[58] = 10'h32b;
        mem[59] = 10'h009;
        mem[60] = 10'h2bc;
        mem[61] = 10'h26b;
        mem[62] = 10'h261;
        mem[63] = 10'h2e1;
        mem[64] = 10'h3db;
        mem[65] = 10'h212;
        mem[66] = 10'h3bd;
        mem[67] = 10'h1ef;
        mem[68] = 10'h229;
        mem[69] = 10'h0c8;
        mem[70] = 10'h187;
        mem[71] = 10'h33d;
        mem[72] = 10'h02e;
        mem[73] = 10'h323;
        mem[74] = 10'h3ce;
        mem[75] = 10'h035;
        mem[76] = 10'h3fa;
        mem[77] = 10'h180;
        mem[78] = 10'h3b9;
        mem[79] = 10'h074;
        mem[80] = 10'h189;
        mem[81] = 10'h372;
        mem[82] = 10'h0a2;
        mem[83] = 10'h383;
        mem[84] = 10'h3b1;
        mem[85] = 10'h207;
        mem[86] = 10'h390;
        mem[87] = 10'h120;
        mem[88] = 10'h30d;
        mem[89] = 10'h33b;
        mem[90] = 10'h001;
        mem[91] = 10'h3ad;
        mem[92] = 10'h391;
        mem[93] = 10'h208;
        mem[94] = 10'h1e6;
        mem[95] = 10'h06e;
        mem[96] = 10'h09f;
        mem[97] = 10'h3cb;
        mem[98] = 10'h2e2;
        mem[99] = 10'h135;
        mem[100] = 10'h3d1;
        mem[101] = 10'h04d;
        mem[102] = 10'h338;
        mem[103] = 10'h0f7;
        mem[104] = 10'h3de;
        mem[105] = 10'h000;
        mem[106] = 10'h317;
        mem[107] = 10'h258;
        mem[108] = 10'h105;
        mem[109] = 10'h1d9;
        mem[110] = 10'h339;
        mem[111] = 10'h24f;
        mem[112] = 10'h289;
        mem[113] = 10'h043;
        mem[114] = 10'h263;
        mem[115] = 10'h332;
        mem[116] = 10'h022;
        mem[117] = 10'h0b6;
        mem[118] = 10'h1ba;
        mem[119] = 10'h098;
        mem[120] = 10'h0ca;
        mem[121] = 10'h1ab;
        mem[122] = 10'h0bf;
        mem[123] = 10'h21b;
        mem[124] = 10'h044;
        mem[125] = 10'h1b7;
        mem[126] = 10'h3b8;
        mem[127] = 10'h3ca;
        mem[128] = 10'h2ee;
        mem[129] = 10'h269;
        mem[130] = 10'h3d9;
        mem[131] = 10'h131;
        mem[132] = 10'h157;
        mem[133] = 10'h089;
        mem[134] = 10'h279;
        mem[135] = 10'h17f;
        mem[136] = 10'h152;
        mem[137] = 10'h25b;
        mem[138] = 10'h214;
        mem[139] = 10'h00e;
        mem[140] = 10'h223;
        mem[141] = 10'h2fd;
        mem[142] = 10'h1dd;
        mem[143] = 10'h199;
        mem[144] = 10'h21d;
        mem[145] = 10'h296;
        mem[146] = 10'h0b4;
        mem[147] = 10'h351;
        mem[148] = 10'h041;
        mem[149] = 10'h03a;
        mem[150] = 10'h201;
        mem[151] = 10'h095;
        mem[152] = 10'h31a;
        mem[153] = 10'h2c0;
        mem[154] = 10'h155;
        mem[155] = 10'h10b;
        mem[156] = 10'h244;
        mem[157] = 10'h1f0;
        mem[158] = 10'h2f7;
        mem[159] = 10'h1f5;
        mem[160] = 10'h227;
        mem[161] = 10'h147;
        mem[162] = 10'h3b6;
        mem[163] = 10'h17c;
        mem[164] = 10'h1c0;
        mem[165] = 10'h094;
        mem[166] = 10'h053;
        mem[167] = 10'h116;
        mem[168] = 10'h245;
        mem[169] = 10'h0dd;
        mem[170] = 10'h2d9;
        mem[171] = 10'h28c;
        mem[172] = 10'h177;
        mem[173] = 10'h3a8;
        mem[174] = 10'h3a4;
        mem[175] = 10'h194;
        mem[176] = 10'h2ce;
        mem[177] = 10'h0ee;
        mem[178] = 10'h172;
        mem[179] = 10'h3f7;
        mem[180] = 10'h0ac;
        mem[181] = 10'h19e;
        mem[182] = 10'h298;
        mem[183] = 10'h134;
        mem[184] = 10'h06f;
        mem[185] = 10'h336;
        mem[186] = 10'h2b8;
        mem[187] = 10'h0dc;
        mem[188] = 10'h33f;
        mem[189] = 10'h05f;
        mem[190] = 10'h1ed;
        mem[191] = 10'h0c9;
        mem[192] = 10'h0ea;
        mem[193] = 10'h1f4;
        mem[194] = 10'h34e;
        mem[195] = 10'h22c;
        mem[196] = 10'h1ad;
        mem[197] = 10'h39c;
        mem[198] = 10'h302;
        mem[199] = 10'h32d;
        mem[200] = 10'h15f;
        mem[201] = 10'h0ef;
        mem[202] = 10'h3fc;
        mem[203] = 10'h108;
        mem[204] = 10'h164;
        mem[205] = 10'h3df;
        mem[206] = 10'h040;
        mem[207] = 10'h084;
        mem[208] = 10'h20b;
        mem[209] = 10'h248;
        mem[210] = 10'h054;
        mem[211] = 10'h0f2;
        mem[212] = 10'h150;
        mem[213] = 10'h01e;
        mem[214] = 10'h11b;
        mem[215] = 10'h2d0;
        mem[216] = 10'h10f;
        mem[217] = 10'h034;
        mem[218] = 10'h3e4;
        mem[219] = 10'h195;
        mem[220] = 10'h38b;
        mem[221] = 10'h119;
        mem[222] = 10'h15c;
        mem[223] = 10'h076;
        mem[224] = 10'h16b;
        mem[225] = 10'h060;
        mem[226] = 10'h114;
        mem[227] = 10'h01d;
        mem[228] = 10'h26c;
        mem[229] = 10'h0da;
        mem[230] = 10'h04e;
        mem[231] = 10'h32e;
        mem[232] = 10'h356;
        mem[233] = 10'h0b3;
        mem[234] = 10'h0c3;
        mem[235] = 10'h1c2;
        mem[236] = 10'h333;
        mem[237] = 10'h253;
        mem[238] = 10'h0e1;
        mem[239] = 10'h3f4;
        mem[240] = 10'h181;
        mem[241] = 10'h14e;
        mem[242] = 10'h20d;
        mem[243] = 10'h138;
        mem[244] = 10'h26e;
        mem[245] = 10'h0c2;
        mem[246] = 10'h15e;
        mem[247] = 10'h216;
        mem[248] = 10'h3cc;
        mem[249] = 10'h3b2;
        mem[250] = 10'h0cc;
        mem[251] = 10'h02c;
        mem[252] = 10'h01f;
        mem[253] = 10'h0c0;
        mem[254] = 10'h230;
        mem[255] = 10'h2a3;
        mem[256] = 10'h2b1;
        mem[257] = 10'h067;
        mem[258] = 10'h1d8;
        mem[259] = 10'h2d2;
        mem[260] = 10'h185;
        mem[261] = 10'h12c;
        mem[262] = 10'h2ea;
        mem[263] = 10'h34f;
        mem[264] = 10'h085;
        mem[265] = 10'h145;
        mem[266] = 10'h0bd;
        mem[267] = 10'h3f9;
        mem[268] = 10'h3a2;
        mem[269] = 10'h0b0;
        mem[270] = 10'h2a4;
        mem[271] = 10'h398;
        mem[272] = 10'h3c6;
        mem[273] = 10'h18f;
        mem[274] = 10'h061;
        mem[275] = 10'h24d;
        mem[276] = 10'h128;
        mem[277] = 10'h273;
        mem[278] = 10'h002;
        mem[279] = 10'h313;
        mem[280] = 10'h2ba;
        mem[281] = 10'h1b9;
        mem[282] = 10'h02d;
        mem[283] = 10'h393;
        mem[284] = 10'h068;
        mem[285] = 10'h361;
        mem[286] = 10'h26a;
        mem[287] = 10'h08c;
        mem[288] = 10'h2c4;
        mem[289] = 10'h109;
        mem[290] = 10'h12d;
        mem[291] = 10'h27d;
        mem[292] = 10'h169;
        mem[293] = 10'h124;
        mem[294] = 10'h047;
        mem[295] = 10'h0f3;
        mem[296] = 10'h10a;
        mem[297] = 10'h3f5;
        mem[298] = 10'h3b5;
        mem[299] = 10'h2d7;
        mem[300] = 10'h02a;
        mem[301] = 10'h0a6;
        mem[302] = 10'h0b5;
        mem[303] = 10'h04c;
        mem[304] = 10'h226;
        mem[305] = 10'h2b3;
        mem[306] = 10'h35f;
        mem[307] = 10'h056;
        mem[308] = 10'h13d;
        mem[309] = 10'h3e9;
        mem[310] = 10'h04a;
        mem[311] = 10'h1f1;
        mem[312] = 10'h2b5;
        mem[313] = 10'h08b;
        mem[314] = 10'h183;
        mem[315] = 10'h06c;
        mem[316] = 10'h17a;
        mem[317] = 10'h0d7;
        mem[318] = 10'h07f;
        mem[319] = 10'h31c;
        mem[320] = 10'h158;
        mem[321] = 10'h295;
        mem[322] = 10'h300;
        mem[323] = 10'h1d0;
        mem[324] = 10'h0f5;
        mem[325] = 10'h0f1;
        mem[326] = 10'h3c4;
        mem[327] = 10'h2ed;
        mem[328] = 10'h274;
        mem[329] = 10'h228;
        mem[330] = 10'h386;
        mem[331] = 10'h003;
        mem[332] = 10'h25a;
        mem[333] = 10'h09d;
        mem[334] = 10'h101;
        mem[335] = 10'h3af;
        mem[336] = 10'h236;
        mem[337] = 10'h1de;
        mem[338] = 10'h104;
        mem[339] = 10'h286;
        mem[340] = 10'h087;
        mem[341] = 10'h0d6;
        mem[342] = 10'h3d6;
        mem[343] = 10'h23a;
        mem[344] = 10'h23c;
        mem[345] = 10'h28e;
        mem[346] = 10'h36f;
        mem[347] = 10'h122;
        mem[348] = 10'h2fb;
        mem[349] = 10'h0f6;
        mem[350] = 10'h3c5;
        mem[351] = 10'h375;
        mem[352] = 10'h11e;
        mem[353] = 10'h1a0;
        mem[354] = 10'h0d8;
        mem[355] = 10'h049;
        mem[356] = 10'h1be;
        mem[357] = 10'h132;
        mem[358] = 10'h112;
        mem[359] = 10'h1b0;
        mem[360] = 10'h051;
        mem[361] = 10'h03c;
        mem[362] = 10'h0a0;
        mem[363] = 10'h00a;
        mem[364] = 10'h384;
        mem[365] = 10'h29e;
        mem[366] = 10'h221;
        mem[367] = 10'h38f;
        mem[368] = 10'h209;
        mem[369] = 10'h357;
        mem[370] = 10'h220;
        mem[371] = 10'h2a5;
        mem[372] = 10'h3d0;
        mem[373] = 10'h37a;
        mem[374] = 10'h345;
        mem[375] = 10'h2e0;
        mem[376] = 10'h0c7;
        mem[377] = 10'h1d2;
        mem[378] = 10'h39e;
        mem[379] = 10'h2e3;
        mem[380] = 10'h26d;
        mem[381] = 10'h280;
        mem[382] = 10'h277;
        mem[383] = 10'h235;
        mem[384] = 10'h2ad;
        mem[385] = 10'h348;
        mem[386] = 10'h0e3;
        mem[387] = 10'h282;
        mem[388] = 10'h048;
        mem[389] = 10'h2e8;
        mem[390] = 10'h330;
        mem[391] = 10'h186;
        mem[392] = 10'h29d;
        mem[393] = 10'h278;
        mem[394] = 10'h34b;
        mem[395] = 10'h005;
        mem[396] = 10'h2e7;
        mem[397] = 10'h373;
        mem[398] = 10'h268;
        mem[399] = 10'h2c3;
        mem[400] = 10'h1ac;
        mem[401] = 10'h1d5;
        mem[402] = 10'h374;
        mem[403] = 10'h2df;
        mem[404] = 10'h0de;
        mem[405] = 10'h140;
        mem[406] = 10'h149;
        mem[407] = 10'h1d7;
        mem[408] = 10'h25c;
        mem[409] = 10'h325;
        mem[410] = 10'h19a;
        mem[411] = 10'h0e7;
        mem[412] = 10'h399;
        mem[413] = 10'h254;
        mem[414] = 10'h2f5;
        mem[415] = 10'h055;
        mem[416] = 10'h0f4;
        mem[417] = 10'h3dd;
        mem[418] = 10'h233;
        mem[419] = 10'h123;
        mem[420] = 10'h1cb;
        mem[421] = 10'h121;
        mem[422] = 10'h246;
        mem[423] = 10'h3c8;
        mem[424] = 10'h340;
        mem[425] = 10'h3e0;
        mem[426] = 10'h0af;
        mem[427] = 10'h163;
        mem[428] = 10'h161;
        mem[429] = 10'h14b;
        mem[430] = 10'h0ff;
        mem[431] = 10'h1ee;
        mem[432] = 10'h1b6;
        mem[433] = 10'h190;
        mem[434] = 10'h030;
        mem[435] = 10'h0fe;
        mem[436] = 10'h35a;
        mem[437] = 10'h3ef;
        mem[438] = 10'h1fb;
        mem[439] = 10'h00c;
        mem[440] = 10'h1da;
        mem[441] = 10'h0e0;
        mem[442] = 10'h24b;
        mem[443] = 10'h362;
        mem[444] = 10'h3be;
        mem[445] = 10'h238;
        mem[446] = 10'h2da;
        mem[447] = 10'h01c;
        mem[448] = 10'h00d;
        mem[449] = 10'h1f9;
        mem[450] = 10'h29c;
        mem[451] = 10'h33c;
        mem[452] = 10'h143;
        mem[453] = 10'h3c7;
        mem[454] = 10'h2ec;
        mem[455] = 10'h275;
        mem[456] = 10'h204;
        mem[457] = 10'h331;
        mem[458] = 10'h2e5;
        mem[459] = 10'h3c1;
        mem[460] = 10'h3e5;
        mem[461] = 10'h0ad;
        mem[462] = 10'h37b;
        mem[463] = 10'h0f0;
        mem[464] = 10'h24c;
        mem[465] = 10'h188;
        mem[466] = 10'h1bc;
        mem[467] = 10'h07c;
        mem[468] = 10'h1e2;
        mem[469] = 10'h290;
        mem[470] = 10'h031;
        mem[471] = 10'h365;
        mem[472] = 10'h14d;
        mem[473] = 10'h3e7;
        mem[474] = 10'h29b;
        mem[475] = 10'h19b;
        mem[476] = 10'h350;
        mem[477] = 10'h353;
        mem[478] = 10'h394;
        mem[479] = 10'h15b;
        mem[480] = 10'h243;
        mem[481] = 10'h37d;
        mem[482] = 10'h100;
        mem[483] = 10'h028;
        mem[484] = 10'h360;
        mem[485] = 10'h2e9;
        mem[486] = 10'h0eb;
        mem[487] = 10'h3aa;
        mem[488] = 10'h262;
        mem[489] = 10'h168;
        mem[490] = 10'h388;
        mem[491] = 10'h08a;
        mem[492] = 10'h3d5;
        mem[493] = 10'h3a6;
        mem[494] = 10'h079;
        mem[495] = 10'h36e;
        mem[496] = 10'h0cf;
        mem[497] = 10'h219;
        mem[498] = 10'h1c4;
        mem[499] = 10'h0b2;
        mem[500] = 10'h2c8;
        mem[501] = 10'h10e;
        mem[502] = 10'h2c1;
        mem[503] = 10'h007;
        mem[504] = 10'h1c5;
        mem[505] = 10'h3a5;
        mem[506] = 10'h2ca;
        mem[507] = 10'h1b1;
        mem[508] = 10'h38e;
        mem[509] = 10'h11d;
        mem[510] = 10'h066;
        mem[511] = 10'h379;
        mem[512] = 10'h1fc;
        mem[513] = 10'h13e;
        mem[514] = 10'h0cb;
        mem[515] = 10'h029;
        mem[516] = 10'h038;
        mem[517] = 10'h0f8;
        mem[518] = 10'h217;
        mem[519] = 10'h04b;
        mem[520] = 10'h255;
        mem[521] = 10'h086;
        mem[522] = 10'h06b;
        mem[523] = 10'h2dd;
        mem[524] = 10'h308;
        mem[525] = 10'h224;
        mem[526] = 10'h0e5;
        mem[527] = 10'h285;
        mem[528] = 10'h242;
        mem[529] = 10'h1c6;
        mem[530] = 10'h1f8;
        mem[531] = 10'h0bc;
        mem[532] = 10'h198;
        mem[533] = 10'h081;
        mem[534] = 10'h0b7;
        mem[535] = 10'h0d2;
        mem[536] = 10'h2b7;
        mem[537] = 10'h213;
        mem[538] = 10'h36d;
        mem[539] = 10'h346;
        mem[540] = 10'h118;
        mem[541] = 10'h320;
        mem[542] = 10'h34d;
        mem[543] = 10'h3bf;
        mem[544] = 10'h0cd;
        mem[545] = 10'h03d;
        mem[546] = 10'h24a;
        mem[547] = 10'h1c1;
        mem[548] = 10'h167;
        mem[549] = 10'h05b;
        mem[550] = 10'h341;
        mem[551] = 10'h3fe;
        mem[552] = 10'h039;
        mem[553] = 10'h178;
        mem[554] = 10'h23b;
        mem[555] = 10'h136;
        mem[556] = 10'h321;
        mem[557] = 10'h1b2;
        mem[558] = 10'h311;
        mem[559] = 10'h3ec;
        mem[560] = 10'h2de;
        mem[561] = 10'h3a7;
        mem[562] = 10'h20c;
        mem[563] = 10'h257;
        mem[564] = 10'h315;
        mem[565] = 10'h385;
        mem[566] = 10'h2d6;
        mem[567] = 10'h160;
        mem[568] = 10'h073;
        mem[569] = 10'h19c;
        mem[570] = 10'h148;
        mem[571] = 10'h1b5;
        mem[572] = 10'h202;
        mem[573] = 10'h04f;
        mem[574] = 10'h1ff;
        mem[575] = 10'h312;
        mem[576] = 10'h2c9;
        mem[577] = 10'h2b0;
        mem[578] = 10'h3b0;
        mem[579] = 10'h144;
        mem[580] = 10'h13b;
        mem[581] = 10'h30c;
        mem[582] = 10'h15a;
        mem[583] = 10'h3cd;
        mem[584] = 10'h106;
        mem[585] = 10'h3f0;
        mem[586] = 10'h111;
        mem[587] = 10'h1a2;
        mem[588] = 10'h21a;
        mem[589] = 10'h1b8;
        mem[590] = 10'h1e1;
        mem[591] = 10'h1ea;
        mem[592] = 10'h17e;
        mem[593] = 10'h03f;
        mem[594] = 10'h082;
        mem[595] = 10'h20e;
        mem[596] = 10'h39f;
        mem[597] = 10'h091;
        mem[598] = 10'h215;
        mem[599] = 10'h32c;
        mem[600] = 10'h03e;
        mem[601] = 10'h39a;
        mem[602] = 10'h058;
        mem[603] = 10'h35e;
        mem[604] = 10'h2a7;
        mem[605] = 10'h080;
        mem[606] = 10'h271;
        mem[607] = 10'h33a;
        mem[608] = 10'h19d;
        mem[609] = 10'h0bb;
        mem[610] = 10'h09b;
        mem[611] = 10'h327;
        mem[612] = 10'h156;
        mem[613] = 10'h283;
        mem[614] = 10'h023;
        mem[615] = 10'h231;
        mem[616] = 10'h1dc;
        mem[617] = 10'h3ee;
        mem[618] = 10'h307;
        mem[619] = 10'h359;
        mem[620] = 10'h267;
        mem[621] = 10'h37c;
        mem[622] = 10'h13c;
        mem[623] = 10'h25f;
        mem[624] = 10'h09c;
        mem[625] = 10'h249;
        mem[626] = 10'h2ef;
        mem[627] = 10'h004;
        mem[628] = 10'h3ff;
        mem[629] = 10'h22f;
        mem[630] = 10'h389;
        mem[631] = 10'h020;
        mem[632] = 10'h38d;
        mem[633] = 10'h162;
        mem[634] = 10'h2bd;
        mem[635] = 10'h2d5;
        mem[636] = 10'h349;
        mem[637] = 10'h059;
        mem[638] = 10'h0ae;
        mem[639] = 10'h3ac;
        mem[640] = 10'h2e4;
        mem[641] = 10'h0fc;
        mem[642] = 10'h38a;
        mem[643] = 10'h057;
        mem[644] = 10'h326;
        mem[645] = 10'h1a5;
        mem[646] = 10'h08d;
        mem[647] = 10'h1ce;
        mem[648] = 10'h09e;
        mem[649] = 10'h09a;
        mem[650] = 10'h3b7;
        mem[651] = 10'h0c1;
        mem[652] = 10'h23e;
        mem[653] = 10'h34c;
        mem[654] = 10'h16a;
        mem[655] = 10'h27a;
        mem[656] = 10'h3d8;
        mem[657] = 10'h011;
        mem[658] = 10'h294;
        mem[659] = 10'h232;
        mem[660] = 10'h0a9;
        mem[661] = 10'h22b;
        mem[662] = 10'h354;
        mem[663] = 10'h166;
        mem[664] = 10'h2d4;
        mem[665] = 10'h0e4;
        mem[666] = 10'h2bb;
        mem[667] = 10'h31b;
        mem[668] = 10'h397;
        mem[669] = 10'h314;
        mem[670] = 10'h026;
        mem[671] = 10'h0be;
        mem[672] = 10'h31d;
        mem[673] = 10'h03b;
        mem[674] = 10'h196;
        mem[675] = 10'h206;
        mem[676] = 10'h130;
        mem[677] = 10'h3ba;
        mem[678] = 10'h069;
        mem[679] = 10'h32f;
        mem[680] = 10'h284;
        mem[681] = 10'h287;
        mem[682] = 10'h033;
        mem[683] = 10'h115;
        mem[684] = 10'h10c;
        mem[685] = 10'h0ab;
        mem[686] = 10'h0b1;
        mem[687] = 10'h0fd;
        mem[688] = 10'h2f0;
        mem[689] = 10'h0a3;
        mem[690] = 10'h26f;
        mem[691] = 10'h304;
        mem[692] = 10'h3e1;
        mem[693] = 10'h0e2;
        mem[694] = 10'h225;
        mem[695] = 10'h38c;
        mem[696] = 10'h20f;
        mem[697] = 10'h133;
        mem[698] = 10'h3d2;
        mem[699] = 10'h1bd;
        mem[700] = 10'h3eb;
        mem[701] = 10'h019;
        mem[702] = 10'h0b8;
        mem[703] = 10'h2ac;
        mem[704] = 10'h0a8;
        mem[705] = 10'h3e6;
        mem[706] = 10'h0d9;
        mem[707] = 10'h1bf;
        mem[708] = 10'h1f6;
        mem[709] = 10'h2cb;
        mem[710] = 10'h1ae;
        mem[711] = 10'h2fa;
        mem[712] = 10'h20a;
        mem[713] = 10'h0ed;
        mem[714] = 10'h16e;
        mem[715] = 10'h259;
        mem[716] = 10'h205;
        mem[717] = 10'h0a4;
        mem[718] = 10'h2cd;
        mem[719] = 10'h3a3;
        mem[720] = 10'h0d5;
        mem[721] = 10'h299;
        mem[722] = 10'h179;
        mem[723] = 10'h088;
        mem[724] = 10'h30e;
        mem[725] = 10'h366;
        mem[726] = 10'h2b6;
        mem[727] = 10'h14a;
        mem[728] = 10'h39b;
        mem[729] = 10'h301;
        mem[730] = 10'h075;
        mem[731] = 10'h2c2;
        mem[732] = 10'h045;
        mem[733] = 10'h1bb;
        mem[734] = 10'h35b;
        mem[735] = 10'h2cf;
        mem[736] = 10'h18c;
        mem[737] = 10'h078;
        mem[738] = 10'h025;
        mem[739] = 10'h3f1;
        mem[740] = 10'h30f;
        mem[741] = 10'h02b;
        mem[742] = 10'h12e;
        mem[743] = 10'h2a0;
        mem[744] = 10'h1cc;
        mem[745] = 10'h2db;
        mem[746] = 10'h309;
        mem[747] = 10'h28a;
        mem[748] = 10'h265;
        mem[749] = 10'h0d0;
        mem[750] = 10'h1e3;
        mem[751] = 10'h395;
        mem[752] = 10'h139;
        mem[753] = 10'h1aa;
        mem[754] = 10'h170;
        mem[755] = 10'h3d7;
        mem[756] = 10'h3ea;
        mem[757] = 10'h305;
        mem[758] = 10'h3ed;
        mem[759] = 10'h050;
        mem[760] = 10'h1c7;
        mem[761] = 10'h18b;
        mem[762] = 10'h16f;
        mem[763] = 10'h2b4;
        mem[764] = 10'h01a;
        mem[765] = 10'h3cf;
        mem[766] = 10'h2f2;
        mem[767] = 10'h1fe;
        mem[768] = 10'h13f;
        mem[769] = 10'h2b2;
        mem[770] = 10'h2c6;
        mem[771] = 10'h18d;
        mem[772] = 10'h381;
        mem[773] = 10'h329;
        mem[774] = 10'h2a8;
        mem[775] = 10'h05d;
        mem[776] = 10'h322;
        mem[777] = 10'h324;
        mem[778] = 10'h2fe;
        mem[779] = 10'h3f3;
        mem[780] = 10'h14c;
        mem[781] = 10'h211;
        mem[782] = 10'h062;
        mem[783] = 10'h16d;
        mem[784] = 10'h200;
        mem[785] = 10'h0ec;
        mem[786] = 10'h376;
        mem[787] = 10'h11a;
        mem[788] = 10'h017;
        mem[789] = 10'h071;
        mem[790] = 10'h08f;
        mem[791] = 10'h103;
        mem[792] = 10'h344;
        mem[793] = 10'h337;
        mem[794] = 10'h264;
        mem[795] = 10'h22e;
        mem[796] = 10'h014;
        mem[797] = 10'h137;
        mem[798] = 10'h1c8;
        mem[799] = 10'h3e3;
        mem[800] = 10'h151;
        mem[801] = 10'h0e9;
        mem[802] = 10'h35d;
        mem[803] = 10'h2bf;
        mem[804] = 10'h1d6;
        mem[805] = 10'h1cf;
        mem[806] = 10'h00f;
        mem[807] = 10'h07a;
        mem[808] = 10'h2f1;
        mem[809] = 10'h016;
        mem[810] = 10'h0d4;
        mem[811] = 10'h024;
        mem[812] = 10'h21f;
        mem[813] = 10'h364;
        mem[814] = 10'h27e;
        mem[815] = 10'h377;
        mem[816] = 10'h21e;
        mem[817] = 10'h1e7;
        mem[818] = 10'h281;
        mem[819] = 10'h127;
        mem[820] = 10'h241;
        mem[821] = 10'h00b;
        mem[822] = 10'h0c5;
        mem[823] = 10'h010;
        mem[824] = 10'h3d4;
        mem[825] = 10'h052;
        mem[826] = 10'h012;
        mem[827] = 10'h29f;
        mem[828] = 10'h36c;
        mem[829] = 10'h27b;
        mem[830] = 10'h032;
        mem[831] = 10'h260;
        mem[832] = 10'h3e2;
        mem[833] = 10'h2d1;
        mem[834] = 10'h102;
        mem[835] = 10'h11c;
        mem[836] = 10'h2c7;
        mem[837] = 10'h15d;
        mem[838] = 10'h318;
        mem[839] = 10'h1d4;
        mem[840] = 10'h070;
        mem[841] = 10'h2f4;
        mem[842] = 10'h07d;
        mem[843] = 10'h0d1;
        mem[844] = 10'h203;
        mem[845] = 10'h256;
        mem[846] = 10'h310;
        mem[847] = 10'h2ae;
        mem[848] = 10'h021;
        mem[849] = 10'h2f9;
        mem[850] = 10'h10d;
        mem[851] = 10'h31f;
        mem[852] = 10'h1fd;
        mem[853] = 10'h008;
        mem[854] = 10'h37e;
        mem[855] = 10'h3e8;
        mem[856] = 10'h0c4;
        mem[857] = 10'h218;
        mem[858] = 10'h25e;
        mem[859] = 10'h083;
        mem[860] = 10'h18a;
        mem[861] = 10'h110;
        mem[862] = 10'h334;
        mem[863] = 10'h3da;
        mem[864] = 10'h1a8;
        mem[865] = 10'h006;
        mem[866] = 10'h065;
        mem[867] = 10'h355;
        mem[868] = 10'h1f7;
        mem[869] = 10'h1e9;
        mem[870] = 10'h342;
        mem[871] = 10'h05a;
        mem[872] = 10'h064;
        mem[873] = 10'h0aa;
        mem[874] = 10'h3bc;
        mem[875] = 10'h2d3;
        mem[876] = 10'h32a;
        mem[877] = 10'h292;
        mem[878] = 10'h1a4;
        mem[879] = 10'h2aa;
        mem[880] = 10'h1e5;
        mem[881] = 10'h1a6;
        mem[882] = 10'h165;
        mem[883] = 10'h0c6;
        mem[884] = 10'h380;
        mem[885] = 10'h2ab;
        mem[886] = 10'h3c9;
        mem[887] = 10'h3c3;
        mem[888] = 10'h37f;
        mem[889] = 10'h2f3;
        mem[890] = 10'h3f6;
        mem[891] = 10'h28b;
        mem[892] = 10'h3dc;
        mem[893] = 10'h3a1;
        mem[894] = 10'h096;
        mem[895] = 10'h18e;
        mem[896] = 10'h015;
        mem[897] = 10'h3f8;
        mem[898] = 10'h01b;
        mem[899] = 10'h293;
        mem[900] = 10'h3ae;
        mem[901] = 10'h23f;
        mem[902] = 10'h3fd;
        mem[903] = 10'h306;
        mem[904] = 10'h22d;
        mem[905] = 10'h247;
        mem[906] = 10'h24e;
        mem[907] = 10'h2cc;
        mem[908] = 10'h358;
        mem[909] = 10'h335;
        mem[910] = 10'h1f2;
        mem[911] = 10'h1a9;
        mem[912] = 10'h1d3;
        mem[913] = 10'h107;
        mem[914] = 10'h018;
        mem[915] = 10'h328;
        mem[916] = 10'h17d;
        mem[917] = 10'h3b3;
        mem[918] = 10'h3b4;
        mem[919] = 10'h1df;
        mem[920] = 10'h34a;
        mem[921] = 10'h0b9;
        mem[922] = 10'h2e6;
        mem[923] = 10'h2f8;
        mem[924] = 10'h382;
        mem[925] = 10'h0ce;
        mem[926] = 10'h1db;
        mem[927] = 10'h240;
        mem[928] = 10'h288;
        mem[929] = 10'h0d3;
        mem[930] = 10'h14f;
        mem[931] = 10'h2d8;
        mem[932] = 10'h171;
        mem[933] = 10'h141;
        mem[934] = 10'h39d;
        mem[935] = 10'h1cd;
        mem[936] = 10'h3a0;
        mem[937] = 10'h22a;
        mem[938] = 10'h1af;
        mem[939] = 10'h35c;
        mem[940] = 10'h2a1;
        mem[941] = 10'h0a1;
        mem[942] = 10'h210;
        mem[943] = 10'h153;
        mem[944] = 10'h30b;
        mem[945] = 10'h36b;
        mem[946] = 10'h396;
        mem[947] = 10'h36a;
        mem[948] = 10'h08e;
        mem[949] = 10'h352;
        mem[950] = 10'h28d;
        mem[951] = 10'h174;
        mem[952] = 10'h129;
        mem[953] = 10'h276;
        mem[954] = 10'h099;
        mem[955] = 10'h042;
        mem[956] = 10'h063;
        mem[957] = 10'h303;
        mem[958] = 10'h251;
        mem[959] = 10'h3f2;
        mem[960] = 10'h05e;
        mem[961] = 10'h270;
        mem[962] = 10'h343;
        mem[963] = 10'h3d3;
        mem[964] = 10'h176;
        mem[965] = 10'h2a6;
        mem[966] = 10'h12a;
        mem[967] = 10'h0df;
        mem[968] = 10'h13a;
        mem[969] = 10'h239;
        mem[970] = 10'h142;
        mem[971] = 10'h192;
        mem[972] = 10'h125;
        mem[973] = 10'h07e;
        mem[974] = 10'h117;
        mem[975] = 10'h072;
        mem[976] = 10'h316;
        mem[977] = 10'h291;
        mem[978] = 10'h21c;
        mem[979] = 10'h2dc;
        mem[980] = 10'h0fb;
        mem[981] = 10'h173;
        mem[982] = 10'h319;
        mem[983] = 10'h1c9;
        mem[984] = 10'h12f;
        mem[985] = 10'h297;
        mem[986] = 10'h17b;
        mem[987] = 10'h154;
        mem[988] = 10'h16c;
        mem[989] = 10'h1fa;
        mem[990] = 10'h387;
        mem[991] = 10'h27c;
        mem[992] = 10'h2f6;
        mem[993] = 10'h27f;
        mem[994] = 10'h12b;
        mem[995] = 10'h146;
        mem[996] = 10'h193;
        mem[997] = 10'h027;
        mem[998] = 10'h06a;
        mem[999] = 10'h0a5;
        mem[1000] = 10'h33e;
        mem[1001] = 10'h28f;
        mem[1002] = 10'h05c;
        mem[1003] = 10'h1a1;
        mem[1004] = 10'h0e6;
        mem[1005] = 10'h378;
        mem[1006] = 10'h1e4;
        mem[1007] = 10'h2fc;
        mem[1008] = 10'h2be;
        mem[1009] = 10'h2af;
        mem[1010] = 10'h1eb;
        mem[1011] = 10'h182;
        mem[1012] = 10'h2a2;
        mem[1013] = 10'h1c3;
        mem[1014] = 10'h0a7;
        mem[1015] = 10'h06d;
        mem[1016] = 10'h184;
        mem[1017] = 10'h369;
        mem[1018] = 10'h3fb;
        mem[1019] = 10'h30a;
        mem[1020] = 10'h1e0;
        mem[1021] = 10'h347;
        mem[1022] = 10'h013;
        mem[1023] = 10'h3a9;
    end
endmodule

module odo_sbox_large5(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    (* ram_style = "block" *) reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h1b9;
        mem[1] = 10'h0ae;
        mem[2] = 10'h2f4;
        mem[3] = 10'h2ed;
        mem[4] = 10'h119;
        mem[5] = 10'h12e;
        mem[6] = 10'h1be;
        mem[7] = 10'h053;
        mem[8] = 10'h349;
        mem[9] = 10'h328;
        mem[10] = 10'h261;
        mem[11] = 10'h24e;
        mem[12] = 10'h06b;
        mem[13] = 10'h165;
        mem[14] = 10'h3f0;
        mem[15] = 10'h249;
        mem[16] = 10'h0af;
        mem[17] = 10'h01c;
        mem[18] = 10'h326;
        mem[19] = 10'h398;
        mem[20] = 10'h21c;
        mem[21] = 10'h3fa;
        mem[22] = 10'h035;
        mem[23] = 10'h32d;
        mem[24] = 10'h05f;
        mem[25] = 10'h00d;
        mem[26] = 10'h108;
        mem[27] = 10'h367;
        mem[28] = 10'h10d;
        mem[29] = 10'h31e;
        mem[30] = 10'h263;
        mem[31] = 10'h259;
        mem[32] = 10'h1d1;
        mem[33] = 10'h106;
        mem[34] = 10'h361;
        mem[35] = 10'h388;
        mem[36] = 10'h015;
        mem[37] = 10'h395;
        mem[38] = 10'h330;
        mem[39] = 10'h3a3;
        mem[40] = 10'h19a;
        mem[41] = 10'h0de;
        mem[42] = 10'h3cc;
        mem[43] = 10'h040;
        mem[44] = 10'h0db;
        mem[45] = 10'h203;
        mem[46] = 10'h1b1;
        mem[47] = 10'h116;
        mem[48] = 10'h3ee;
        mem[49] = 10'h22e;
        mem[50] = 10'h3b8;
        mem[51] = 10'h064;
        mem[52] = 10'h0fb;
        mem[53] = 10'h1a3;
        mem[54] = 10'h0ab;
        mem[55] = 10'h3b2;
        mem[56] = 10'h2c8;
        mem[57] = 10'h375;
        mem[58] = 10'h078;
        mem[59] = 10'h1d2;
        mem[60] = 10'h074;
        mem[61] = 10'h317;
        mem[62] = 10'h009;
        mem[63] = 10'h00e;
        mem[64] = 10'h000;
        mem[65] = 10'h32a;
        mem[66] = 10'h1eb;
        mem[67] = 10'h08b;
        mem[68] = 10'h2ec;
        mem[69] = 10'h3a1;
        mem[70] = 10'h312;
        mem[71] = 10'h1ed;
        mem[72] = 10'h2d9;
        mem[73] = 10'h39e;
        mem[74] = 10'h1ea;
        mem[75] = 10'h0b3;
        mem[76] = 10'h20b;
        mem[77] = 10'h122;
        mem[78] = 10'h077;
        mem[79] = 10'h120;
        mem[80] = 10'h05c;
        mem[81] = 10'h189;
        mem[82] = 10'h1df;
        mem[83] = 10'h05d;
        mem[84] = 10'h0d9;
        mem[85] = 10'h002;
        mem[86] = 10'h18b;
        mem[87] = 10'h0d4;
        mem[88] = 10'h012;
        mem[89] = 10'h0c2;
        mem[90] = 10'h3db;
        mem[91] = 10'h3f8;
        mem[92] = 10'h223;
        mem[93] = 10'h31f;
        mem[94] = 10'h030;
        mem[95] = 10'h2b9;
        mem[96] = 10'h284;
        mem[97] = 10'h04a;
        mem[98] = 10'h3e3;
        mem[99] = 10'h2b0;
        mem[100] = 10'h10b;
        mem[101] = 10'h258;
        mem[102] = 10'h1d5;
        mem[103] = 10'h228;
        mem[104] = 10'h2a9;
        mem[105] = 10'h07c;
        mem[106] = 10'h368;
        mem[107] = 10'h117;
        mem[108] = 10'h16b;
        mem[109] = 10'h260;
        mem[110] = 10'h0c1;
        mem[111] = 10'h3cd;
        mem[112] = 10'h36a;
        mem[113] = 10'h147;
        mem[114] = 10'h07a;
        mem[115] = 10'h1da;
        mem[116] = 10'h0ce;
        mem[117] = 10'h3a9;
        mem[118] = 10'h335;
        mem[119] = 10'h156;
        mem[120] = 10'h1f8;
        mem[121] = 10'h073;
        mem[122] = 10'h2a1;
        mem[123] = 10'h220;
        mem[124] = 10'h33e;
        mem[125] = 10'h101;
        mem[126] = 10'h36d;
        mem[127] = 10'h288;
        mem[128] = 10'h3d0;
        mem[129] = 10'h2cd;
        mem[130] = 10'h344;
        mem[131] = 10'h313;
        mem[132] = 10'h10e;
        mem[133] = 10'h01e;
        mem[134] = 10'h38a;
        mem[135] = 10'h3ae;
        mem[136] = 10'h3d4;
        mem[137] = 10'h04d;
        mem[138] = 10'h121;
        mem[139] = 10'h18f;
        mem[140] = 10'h3f2;
        mem[141] = 10'h0a0;
        mem[142] = 10'h25b;
        mem[143] = 10'h2cf;
        mem[144] = 10'h0bb;
        mem[145] = 10'h378;
        mem[146] = 10'h216;
        mem[147] = 10'h1c6;
        mem[148] = 10'h204;
        mem[149] = 10'h3a7;
        mem[150] = 10'h3aa;
        mem[151] = 10'h327;
        mem[152] = 10'h294;
        mem[153] = 10'h227;
        mem[154] = 10'h018;
        mem[155] = 10'h23f;
        mem[156] = 10'h1d4;
        mem[157] = 10'h24b;
        mem[158] = 10'h16d;
        mem[159] = 10'h27d;
        mem[160] = 10'h148;
        mem[161] = 10'h0b0;
        mem[162] = 10'h177;
        mem[163] = 10'h04b;
        mem[164] = 10'h353;
        mem[165] = 10'h039;
        mem[166] = 10'h2fa;
        mem[167] = 10'h2cc;
        mem[168] = 10'h303;
        mem[169] = 10'h180;
        mem[170] = 10'h379;
        mem[171] = 10'h098;
        mem[172] = 10'h345;
        mem[173] = 10'h38c;
        mem[174] = 10'h0e8;
        mem[175] = 10'h214;
        mem[176] = 10'h16a;
        mem[177] = 10'h09c;
        mem[178] = 10'h0bc;
        mem[179] = 10'h221;
        mem[180] = 10'h2e8;
        mem[181] = 10'h371;
        mem[182] = 10'h1c1;
        mem[183] = 10'h05b;
        mem[184] = 10'h2a4;
        mem[185] = 10'h26b;
        mem[186] = 10'h022;
        mem[187] = 10'h01b;
        mem[188] = 10'h065;
        mem[189] = 10'h0f5;
        mem[190] = 10'h3c6;
        mem[191] = 10'h10c;
        mem[192] = 10'h332;
        mem[193] = 10'h369;
        mem[194] = 10'h280;
        mem[195] = 10'h113;
        mem[196] = 10'h1d8;
        mem[197] = 10'h0b2;
        mem[198] = 10'h070;
        mem[199] = 10'h22c;
        mem[200] = 10'h295;
        mem[201] = 10'h231;
        mem[202] = 10'h0e3;
        mem[203] = 10'h36f;
        mem[204] = 10'h20e;
        mem[205] = 10'h055;
        mem[206] = 10'h096;
        mem[207] = 10'h004;
        mem[208] = 10'h318;
        mem[209] = 10'h338;
        mem[210] = 10'h03a;
        mem[211] = 10'h083;
        mem[212] = 10'h3d5;
        mem[213] = 10'h2ff;
        mem[214] = 10'h19d;
        mem[215] = 10'h2c4;
        mem[216] = 10'h2b1;
        mem[217] = 10'h26c;
        mem[218] = 10'h010;
        mem[219] = 10'h182;
        mem[220] = 10'h0cd;
        mem[221] = 10'h3dc;
        mem[222] = 10'h244;
        mem[223] = 10'h0a4;
        mem[224] = 10'h1b6;
        mem[225] = 10'h18d;
        mem[226] = 10'h136;
        mem[227] = 10'h2b3;
        mem[228] = 10'h0a3;
        mem[229] = 10'h38d;
        mem[230] = 10'h289;
        mem[231] = 10'h008;
        mem[232] = 10'h28b;
        mem[233] = 10'h157;
        mem[234] = 10'h179;
        mem[235] = 10'h050;
        mem[236] = 10'h2f5;
        mem[237] = 10'h22d;
        mem[238] = 10'h27a;
        mem[239] = 10'h15a;
        mem[240] = 10'h274;
        mem[241] = 10'h1a9;
        mem[242] = 10'h1dd;
        mem[243] = 10'h381;
        mem[244] = 10'h391;
        mem[245] = 10'h3e0;
        mem[246] = 10'h08f;
        mem[247] = 10'h287;
        mem[248] = 10'h187;
        mem[249] = 10'h115;
        mem[250] = 10'h28f;
        mem[251] = 10'h13d;
        mem[252] = 10'h1e2;
        mem[253] = 10'h3f1;
        mem[254] = 10'h0b7;
        mem[255] = 10'h30f;
        mem[256] = 10'h2fb;
        mem[257] = 10'h1bc;
        mem[258] = 10'h2df;
        mem[259] = 10'h2b8;
        mem[260] = 10'h235;
        mem[261] = 10'h105;
        mem[262] = 10'h128;
        mem[263] = 10'h2f1;
        mem[264] = 10'h3a5;
        mem[265] = 10'h14f;
        mem[266] = 10'h2fe;
        mem[267] = 10'h333;
        mem[268] = 10'h123;
        mem[269] = 10'h019;
        mem[270] = 10'h1fc;
        mem[271] = 10'h201;
        mem[272] = 10'h269;
        mem[273] = 10'h14b;
        mem[274] = 10'h18a;
        mem[275] = 10'h270;
        mem[276] = 10'h2a5;
        mem[277] = 10'h256;
        mem[278] = 10'h06d;
        mem[279] = 10'h153;
        mem[280] = 10'h2a0;
        mem[281] = 10'h250;
        mem[282] = 10'h3d6;
        mem[283] = 10'h0c5;
        mem[284] = 10'h320;
        mem[285] = 10'h2c7;
        mem[286] = 10'h2c1;
        mem[287] = 10'h2e6;
        mem[288] = 10'h152;
        mem[289] = 10'h141;
        mem[290] = 10'h307;
        mem[291] = 10'h217;
        mem[292] = 10'h208;
        mem[293] = 10'h3c2;
        mem[294] = 10'h296;
        mem[295] = 10'h308;
        mem[296] = 10'h35a;
        mem[297] = 10'h03e;
        mem[298] = 10'h255;
        mem[299] = 10'h170;
        mem[300] = 10'h253;
        mem[301] = 10'h13c;
        mem[302] = 10'h3ba;
        mem[303] = 10'h1a2;
        mem[304] = 10'h215;
        mem[305] = 10'h0c8;
        mem[306] = 10'h2b6;
        mem[307] = 10'h0e6;
        mem[308] = 10'h1af;
        mem[309] = 10'h1c0;
        mem[310] = 10'h0a8;
        mem[311] = 10'h134;
        mem[312] = 10'h3bc;
        mem[313] = 10'h3c1;
        mem[314] = 10'h1b7;
        mem[315] = 10'h20a;
        mem[316] = 10'h362;
        mem[317] = 10'h049;
        mem[318] = 10'h315;
        mem[319] = 10'h02c;
        mem[320] = 10'h241;
        mem[321] = 10'h0f3;
        mem[322] = 10'h0ed;
        mem[323] = 10'h310;
        mem[324] = 10'h396;
        mem[325] = 10'h286;
        mem[326] = 10'h3ec;
        mem[327] = 10'h17b;
        mem[328] = 10'h202;
        mem[329] = 10'h384;
        mem[330] = 10'h192;
        mem[331] = 10'h0be;
        mem[332] = 10'h06c;
        mem[333] = 10'h20c;
        mem[334] = 10'h033;
        mem[335] = 10'h185;
        mem[336] = 10'h33a;
        mem[337] = 10'h370;
        mem[338] = 10'h27e;
        mem[339] = 10'h211;
        mem[340] = 10'h3eb;
        mem[341] = 10'h09f;
        mem[342] = 10'h278;
        mem[343] = 10'h32e;
        mem[344] = 10'h11f;
        mem[345] = 10'h2ce;
        mem[346] = 10'h0f0;
        mem[347] = 10'h1e4;
        mem[348] = 10'h042;
        mem[349] = 10'h100;
        mem[350] = 10'h10a;
        mem[351] = 10'h373;
        mem[352] = 10'h2f0;
        mem[353] = 10'h162;
        mem[354] = 10'h3d2;
        mem[355] = 10'h2de;
        mem[356] = 10'h0eb;
        mem[357] = 10'h277;
        mem[358] = 10'h2f3;
        mem[359] = 10'h005;
        mem[360] = 10'h14c;
        mem[361] = 10'h27f;
        mem[362] = 10'h3e9;
        mem[363] = 10'h37d;
        mem[364] = 10'h1d7;
        mem[365] = 10'h1a5;
        mem[366] = 10'h158;
        mem[367] = 10'h2ac;
        mem[368] = 10'h299;
        mem[369] = 10'h107;
        mem[370] = 10'h087;
        mem[371] = 10'h32f;
        mem[372] = 10'h268;
        mem[373] = 10'h2a8;
        mem[374] = 10'h390;
        mem[375] = 10'h23d;
        mem[376] = 10'h1fa;
        mem[377] = 10'h020;
        mem[378] = 10'h266;
        mem[379] = 10'h397;
        mem[380] = 10'h16f;
        mem[381] = 10'h3ed;
        mem[382] = 10'h2bc;
        mem[383] = 10'h2e1;
        mem[384] = 10'h39c;
        mem[385] = 10'h2f8;
        mem[386] = 10'h350;
        mem[387] = 10'h00f;
        mem[388] = 10'h0a9;
        mem[389] = 10'h355;
        mem[390] = 10'h043;
        mem[391] = 10'h1ff;
        mem[392] = 10'h2d8;
        mem[393] = 10'h0d7;
        mem[394] = 10'h285;
        mem[395] = 10'h0e1;
        mem[396] = 10'h324;
        mem[397] = 10'h2b2;
        mem[398] = 10'h264;
        mem[399] = 10'h12a;
        mem[400] = 10'h02f;
        mem[401] = 10'h321;
        mem[402] = 10'h1f6;
        mem[403] = 10'h3a0;
        mem[404] = 10'h3dd;
        mem[405] = 10'h3be;
        mem[406] = 10'h1cb;
        mem[407] = 10'h026;
        mem[408] = 10'h17f;
        mem[409] = 10'h1ce;
        mem[410] = 10'h3c9;
        mem[411] = 10'h17c;
        mem[412] = 10'h316;
        mem[413] = 10'h0d1;
        mem[414] = 10'h267;
        mem[415] = 10'h3f7;
        mem[416] = 10'h305;
        mem[417] = 10'h173;
        mem[418] = 10'h1ba;
        mem[419] = 10'h314;
        mem[420] = 10'h1ca;
        mem[421] = 10'h2b4;
        mem[422] = 10'h06f;
        mem[423] = 10'h13e;
        mem[424] = 10'h209;
        mem[425] = 10'h1e8;
        mem[426] = 10'h1a1;
        mem[427] = 10'h054;
        mem[428] = 10'h240;
        mem[429] = 10'h021;
        mem[430] = 10'h1de;
        mem[431] = 10'h178;
        mem[432] = 10'h32b;
        mem[433] = 10'h144;
        mem[434] = 10'h357;
        mem[435] = 10'h079;
        mem[436] = 10'h1fd;
        mem[437] = 10'h26f;
        mem[438] = 10'h2a6;
        mem[439] = 10'h19e;
        mem[440] = 10'h239;
        mem[441] = 10'h3fc;
        mem[442] = 10'h02e;
        mem[443] = 10'h1b0;
        mem[444] = 10'h2c6;
        mem[445] = 10'h3af;
        mem[446] = 10'h032;
        mem[447] = 10'h12d;
        mem[448] = 10'h3c4;
        mem[449] = 10'h15f;
        mem[450] = 10'h155;
        mem[451] = 10'h1ee;
        mem[452] = 10'h3cf;
        mem[453] = 10'h34e;
        mem[454] = 10'h218;
        mem[455] = 10'h2e9;
        mem[456] = 10'h257;
        mem[457] = 10'h2ba;
        mem[458] = 10'h243;
        mem[459] = 10'h0ea;
        mem[460] = 10'h392;
        mem[461] = 10'h1bd;
        mem[462] = 10'h2ab;
        mem[463] = 10'h3a6;
        mem[464] = 10'h2e5;
        mem[465] = 10'h011;
        mem[466] = 10'h052;
        mem[467] = 10'h0b4;
        mem[468] = 10'h15e;
        mem[469] = 10'h3b4;
        mem[470] = 10'h29e;
        mem[471] = 10'h2be;
        mem[472] = 10'h1c9;
        mem[473] = 10'h279;
        mem[474] = 10'h02d;
        mem[475] = 10'h1c3;
        mem[476] = 10'h36b;
        mem[477] = 10'h339;
        mem[478] = 10'h23e;
        mem[479] = 10'h061;
        mem[480] = 10'h376;
        mem[481] = 10'h33f;
        mem[482] = 10'h325;
        mem[483] = 10'h394;
        mem[484] = 10'h034;
        mem[485] = 10'h07d;
        mem[486] = 10'h1a0;
        mem[487] = 10'h38e;
        mem[488] = 10'h2d0;
        mem[489] = 10'h0b8;
        mem[490] = 10'h03b;
        mem[491] = 10'h348;
        mem[492] = 10'h03d;
        mem[493] = 10'h31c;
        mem[494] = 10'h071;
        mem[495] = 10'h275;
        mem[496] = 10'h2bf;
        mem[497] = 10'h14d;
        mem[498] = 10'h198;
        mem[499] = 10'h200;
        mem[500] = 10'h232;
        mem[501] = 10'h3b7;
        mem[502] = 10'h0cb;
        mem[503] = 10'h38f;
        mem[504] = 10'h30b;
        mem[505] = 10'h340;
        mem[506] = 10'h0aa;
        mem[507] = 10'h090;
        mem[508] = 10'h283;
        mem[509] = 10'h031;
        mem[510] = 10'h12c;
        mem[511] = 10'h013;
        mem[512] = 10'h11b;
        mem[513] = 10'h10f;
        mem[514] = 10'h0c3;
        mem[515] = 10'h150;
        mem[516] = 10'h1f0;
        mem[517] = 10'h3ab;
        mem[518] = 10'h139;
        mem[519] = 10'h29d;
        mem[520] = 10'h2c3;
        mem[521] = 10'h1e0;
        mem[522] = 10'h251;
        mem[523] = 10'h2da;
        mem[524] = 10'h15c;
        mem[525] = 10'h159;
        mem[526] = 10'h293;
        mem[527] = 10'h0b5;
        mem[528] = 10'h06e;
        mem[529] = 10'h27c;
        mem[530] = 10'h1d3;
        mem[531] = 10'h23b;
        mem[532] = 10'h1e7;
        mem[533] = 10'h230;
        mem[534] = 10'h048;
        mem[535] = 10'h358;
        mem[536] = 10'h3f9;
        mem[537] = 10'h21a;
        mem[538] = 10'h21b;
        mem[539] = 10'h0a5;
        mem[540] = 10'h3f3;
        mem[541] = 10'h309;
        mem[542] = 10'h298;
        mem[543] = 10'h3e8;
        mem[544] = 10'h1fb;
        mem[545] = 10'h39b;
        mem[546] = 10'h023;
        mem[547] = 10'h35e;
        mem[548] = 10'h245;
        mem[549] = 10'h302;
        mem[550] = 10'h0a1;
        mem[551] = 10'h2a3;
        mem[552] = 10'h0f6;
        mem[553] = 10'h0e7;
        mem[554] = 10'h2d5;
        mem[555] = 10'h20f;
        mem[556] = 10'h399;
        mem[557] = 10'h1f7;
        mem[558] = 10'h114;
        mem[559] = 10'h39f;
        mem[560] = 10'h11c;
        mem[561] = 10'h0b6;
        mem[562] = 10'h0b9;
        mem[563] = 10'h2af;
        mem[564] = 10'h069;
        mem[565] = 10'h197;
        mem[566] = 10'h0e9;
        mem[567] = 10'h25c;
        mem[568] = 10'h304;
        mem[569] = 10'h2ae;
        mem[570] = 10'h2c9;
        mem[571] = 10'h2e7;
        mem[572] = 10'h25a;
        mem[573] = 10'h39a;
        mem[574] = 10'h1ab;
        mem[575] = 10'h290;
        mem[576] = 10'h3ac;
        mem[577] = 10'h380;
        mem[578] = 10'h140;
        mem[579] = 10'h2bd;
        mem[580] = 10'h137;
        mem[581] = 10'h0d0;
        mem[582] = 10'h2b7;
        mem[583] = 10'h01a;
        mem[584] = 10'h095;
        mem[585] = 10'h364;
        mem[586] = 10'h347;
        mem[587] = 10'h01d;
        mem[588] = 10'h36c;
        mem[589] = 10'h14a;
        mem[590] = 10'h1f2;
        mem[591] = 10'h24c;
        mem[592] = 10'h354;
        mem[593] = 10'h169;
        mem[594] = 10'h246;
        mem[595] = 10'h027;
        mem[596] = 10'h24a;
        mem[597] = 10'h3b0;
        mem[598] = 10'h3b6;
        mem[599] = 10'h068;
        mem[600] = 10'h219;
        mem[601] = 10'h13f;
        mem[602] = 10'h19c;
        mem[603] = 10'h33c;
        mem[604] = 10'h3c0;
        mem[605] = 10'h082;
        mem[606] = 10'h3a2;
        mem[607] = 10'h3ef;
        mem[608] = 10'h024;
        mem[609] = 10'h199;
        mem[610] = 10'h1c7;
        mem[611] = 10'h03c;
        mem[612] = 10'h0d5;
        mem[613] = 10'h3d7;
        mem[614] = 10'h176;
        mem[615] = 10'h3cb;
        mem[616] = 10'h01f;
        mem[617] = 10'h0a7;
        mem[618] = 10'h1dc;
        mem[619] = 10'h196;
        mem[620] = 10'h3c7;
        mem[621] = 10'h3c5;
        mem[622] = 10'h058;
        mem[623] = 10'h2d3;
        mem[624] = 10'h02a;
        mem[625] = 10'h051;
        mem[626] = 10'h184;
        mem[627] = 10'h3b3;
        mem[628] = 10'h190;
        mem[629] = 10'h22b;
        mem[630] = 10'h0ee;
        mem[631] = 10'h14e;
        mem[632] = 10'h036;
        mem[633] = 10'h236;
        mem[634] = 10'h0dc;
        mem[635] = 10'h3e7;
        mem[636] = 10'h191;
        mem[637] = 10'h25e;
        mem[638] = 10'h142;
        mem[639] = 10'h30d;
        mem[640] = 10'h31a;
        mem[641] = 10'h04f;
        mem[642] = 10'h18c;
        mem[643] = 10'h19f;
        mem[644] = 10'h08c;
        mem[645] = 10'h126;
        mem[646] = 10'h1d6;
        mem[647] = 10'h0bd;
        mem[648] = 10'h2dd;
        mem[649] = 10'h24d;
        mem[650] = 10'h276;
        mem[651] = 10'h047;
        mem[652] = 10'h2c0;
        mem[653] = 10'h112;
        mem[654] = 10'h00b;
        mem[655] = 10'h138;
        mem[656] = 10'h21e;
        mem[657] = 10'h3ca;
        mem[658] = 10'h081;
        mem[659] = 10'h3fd;
        mem[660] = 10'h1ad;
        mem[661] = 10'h11a;
        mem[662] = 10'h33b;
        mem[663] = 10'h1a6;
        mem[664] = 10'h1e9;
        mem[665] = 10'h09e;
        mem[666] = 10'h0ca;
        mem[667] = 10'h08d;
        mem[668] = 10'h067;
        mem[669] = 10'h086;
        mem[670] = 10'h2f6;
        mem[671] = 10'h017;
        mem[672] = 10'h102;
        mem[673] = 10'h181;
        mem[674] = 10'h0fc;
        mem[675] = 10'h20d;
        mem[676] = 10'h161;
        mem[677] = 10'h066;
        mem[678] = 10'h34c;
        mem[679] = 10'h366;
        mem[680] = 10'h2b5;
        mem[681] = 10'h038;
        mem[682] = 10'h063;
        mem[683] = 10'h3e5;
        mem[684] = 10'h3df;
        mem[685] = 10'h0a6;
        mem[686] = 10'h3b9;
        mem[687] = 10'h2eb;
        mem[688] = 10'h30c;
        mem[689] = 10'h103;
        mem[690] = 10'h1ec;
        mem[691] = 10'h2d7;
        mem[692] = 10'h014;
        mem[693] = 10'h21f;
        mem[694] = 10'h3bf;
        mem[695] = 10'h252;
        mem[696] = 10'h154;
        mem[697] = 10'h3fe;
        mem[698] = 10'h0f8;
        mem[699] = 10'h301;
        mem[700] = 10'h1bb;
        mem[701] = 10'h300;
        mem[702] = 10'h0ef;
        mem[703] = 10'h206;
        mem[704] = 10'h05a;
        mem[705] = 10'h016;
        mem[706] = 10'h075;
        mem[707] = 10'h124;
        mem[708] = 10'h291;
        mem[709] = 10'h2a7;
        mem[710] = 10'h127;
        mem[711] = 10'h32c;
        mem[712] = 10'h29b;
        mem[713] = 10'h319;
        mem[714] = 10'h072;
        mem[715] = 10'h272;
        mem[716] = 10'h17d;
        mem[717] = 10'h30a;
        mem[718] = 10'h1b5;
        mem[719] = 10'h045;
        mem[720] = 10'h092;
        mem[721] = 10'h12b;
        mem[722] = 10'h3f5;
        mem[723] = 10'h125;
        mem[724] = 10'h046;
        mem[725] = 10'h35c;
        mem[726] = 10'h28a;
        mem[727] = 10'h323;
        mem[728] = 10'h060;
        mem[729] = 10'h2f7;
        mem[730] = 10'h3e6;
        mem[731] = 10'h242;
        mem[732] = 10'h135;
        mem[733] = 10'h149;
        mem[734] = 10'h0d8;
        mem[735] = 10'h171;
        mem[736] = 10'h1b2;
        mem[737] = 10'h3da;
        mem[738] = 10'h234;
        mem[739] = 10'h37e;
        mem[740] = 10'h110;
        mem[741] = 10'h39d;
        mem[742] = 10'h00c;
        mem[743] = 10'h359;
        mem[744] = 10'h0d3;
        mem[745] = 10'h3d3;
        mem[746] = 10'h09a;
        mem[747] = 10'h386;
        mem[748] = 10'h0ad;
        mem[749] = 10'h374;
        mem[750] = 10'h1a7;
        mem[751] = 10'h282;
        mem[752] = 10'h194;
        mem[753] = 10'h1c2;
        mem[754] = 10'h2e3;
        mem[755] = 10'h1aa;
        mem[756] = 10'h22a;
        mem[757] = 10'h372;
        mem[758] = 10'h037;
        mem[759] = 10'h15d;
        mem[760] = 10'h336;
        mem[761] = 10'h352;
        mem[762] = 10'h37f;
        mem[763] = 10'h168;
        mem[764] = 10'h205;
        mem[765] = 10'h3c8;
        mem[766] = 10'h0f1;
        mem[767] = 10'h1d9;
        mem[768] = 10'h2ad;
        mem[769] = 10'h334;
        mem[770] = 10'h3fb;
        mem[771] = 10'h3f4;
        mem[772] = 10'h238;
        mem[773] = 10'h226;
        mem[774] = 10'h1e5;
        mem[775] = 10'h233;
        mem[776] = 10'h08a;
        mem[777] = 10'h059;
        mem[778] = 10'h363;
        mem[779] = 10'h146;
        mem[780] = 10'h1b8;
        mem[781] = 10'h1f5;
        mem[782] = 10'h05e;
        mem[783] = 10'h1b4;
        mem[784] = 10'h0c7;
        mem[785] = 10'h097;
        mem[786] = 10'h0e4;
        mem[787] = 10'h1a8;
        mem[788] = 10'h1e6;
        mem[789] = 10'h1f4;
        mem[790] = 10'h29f;
        mem[791] = 10'h262;
        mem[792] = 10'h329;
        mem[793] = 10'h025;
        mem[794] = 10'h172;
        mem[795] = 10'h2d4;
        mem[796] = 10'h2d2;
        mem[797] = 10'h00a;
        mem[798] = 10'h2c2;
        mem[799] = 10'h3ff;
        mem[800] = 10'h1ac;
        mem[801] = 10'h31b;
        mem[802] = 10'h3e2;
        mem[803] = 10'h09d;
        mem[804] = 10'h2cb;
        mem[805] = 10'h2ee;
        mem[806] = 10'h3d8;
        mem[807] = 10'h001;
        mem[808] = 10'h044;
        mem[809] = 10'h2f2;
        mem[810] = 10'h13b;
        mem[811] = 10'h254;
        mem[812] = 10'h174;
        mem[813] = 10'h104;
        mem[814] = 10'h34a;
        mem[815] = 10'h085;
        mem[816] = 10'h281;
        mem[817] = 10'h207;
        mem[818] = 10'h0fd;
        mem[819] = 10'h163;
        mem[820] = 10'h16e;
        mem[821] = 10'h311;
        mem[822] = 10'h007;
        mem[823] = 10'h34f;
        mem[824] = 10'h151;
        mem[825] = 10'h0bf;
        mem[826] = 10'h0ba;
        mem[827] = 10'h1e1;
        mem[828] = 10'h385;
        mem[829] = 10'h2aa;
        mem[830] = 10'h29a;
        mem[831] = 10'h17e;
        mem[832] = 10'h351;
        mem[833] = 10'h0df;
        mem[834] = 10'h31d;
        mem[835] = 10'h360;
        mem[836] = 10'h1cf;
        mem[837] = 10'h387;
        mem[838] = 10'h0c6;
        mem[839] = 10'h0fe;
        mem[840] = 10'h080;
        mem[841] = 10'h2ca;
        mem[842] = 10'h346;
        mem[843] = 10'h143;
        mem[844] = 10'h331;
        mem[845] = 10'h3bd;
        mem[846] = 10'h365;
        mem[847] = 10'h2fc;
        mem[848] = 10'h2e4;
        mem[849] = 10'h1c4;
        mem[850] = 10'h389;
        mem[851] = 10'h1ae;
        mem[852] = 10'h0c9;
        mem[853] = 10'h076;
        mem[854] = 10'h306;
        mem[855] = 10'h094;
        mem[856] = 10'h188;
        mem[857] = 10'h13a;
        mem[858] = 10'h028;
        mem[859] = 10'h28e;
        mem[860] = 10'h393;
        mem[861] = 10'h11d;
        mem[862] = 10'h229;
        mem[863] = 10'h2c5;
        mem[864] = 10'h3a8;
        mem[865] = 10'h0f9;
        mem[866] = 10'h225;
        mem[867] = 10'h3a4;
        mem[868] = 10'h3e1;
        mem[869] = 10'h2f9;
        mem[870] = 10'h0f2;
        mem[871] = 10'h222;
        mem[872] = 10'h3bb;
        mem[873] = 10'h356;
        mem[874] = 10'h382;
        mem[875] = 10'h16c;
        mem[876] = 10'h35b;
        mem[877] = 10'h271;
        mem[878] = 10'h224;
        mem[879] = 10'h08e;
        mem[880] = 10'h3b5;
        mem[881] = 10'h118;
        mem[882] = 10'h041;
        mem[883] = 10'h006;
        mem[884] = 10'h04c;
        mem[885] = 10'h2ea;
        mem[886] = 10'h133;
        mem[887] = 10'h129;
        mem[888] = 10'h130;
        mem[889] = 10'h1d0;
        mem[890] = 10'h3de;
        mem[891] = 10'h37b;
        mem[892] = 10'h2a2;
        mem[893] = 10'h003;
        mem[894] = 10'h297;
        mem[895] = 10'h195;
        mem[896] = 10'h1c5;
        mem[897] = 10'h164;
        mem[898] = 10'h07f;
        mem[899] = 10'h1c8;
        mem[900] = 10'h0a2;
        mem[901] = 10'h26e;
        mem[902] = 10'h2d1;
        mem[903] = 10'h07b;
        mem[904] = 10'h3d1;
        mem[905] = 10'h337;
        mem[906] = 10'h17a;
        mem[907] = 10'h0ac;
        mem[908] = 10'h35f;
        mem[909] = 10'h30e;
        mem[910] = 10'h292;
        mem[911] = 10'h2d6;
        mem[912] = 10'h0b1;
        mem[913] = 10'h2fd;
        mem[914] = 10'h21d;
        mem[915] = 10'h0e0;
        mem[916] = 10'h34b;
        mem[917] = 10'h091;
        mem[918] = 10'h0fa;
        mem[919] = 10'h3d9;
        mem[920] = 10'h193;
        mem[921] = 10'h3c3;
        mem[922] = 10'h2e0;
        mem[923] = 10'h145;
        mem[924] = 10'h0da;
        mem[925] = 10'h12f;
        mem[926] = 10'h25d;
        mem[927] = 10'h2e2;
        mem[928] = 10'h04e;
        mem[929] = 10'h07e;
        mem[930] = 10'h23c;
        mem[931] = 10'h3e4;
        mem[932] = 10'h0cc;
        mem[933] = 10'h37c;
        mem[934] = 10'h2db;
        mem[935] = 10'h0d6;
        mem[936] = 10'h3f6;
        mem[937] = 10'h322;
        mem[938] = 10'h09b;
        mem[939] = 10'h06a;
        mem[940] = 10'h343;
        mem[941] = 10'h212;
        mem[942] = 10'h062;
        mem[943] = 10'h0dd;
        mem[944] = 10'h183;
        mem[945] = 10'h210;
        mem[946] = 10'h166;
        mem[947] = 10'h175;
        mem[948] = 10'h3ea;
        mem[949] = 10'h29c;
        mem[950] = 10'h1cc;
        mem[951] = 10'h2ef;
        mem[952] = 10'h099;
        mem[953] = 10'h056;
        mem[954] = 10'h1b3;
        mem[955] = 10'h03f;
        mem[956] = 10'h1ef;
        mem[957] = 10'h131;
        mem[958] = 10'h084;
        mem[959] = 10'h1f9;
        mem[960] = 10'h160;
        mem[961] = 10'h3ce;
        mem[962] = 10'h0e5;
        mem[963] = 10'h342;
        mem[964] = 10'h093;
        mem[965] = 10'h186;
        mem[966] = 10'h1f1;
        mem[967] = 10'h089;
        mem[968] = 10'h27b;
        mem[969] = 10'h132;
        mem[970] = 10'h0d2;
        mem[971] = 10'h28c;
        mem[972] = 10'h18e;
        mem[973] = 10'h1f3;
        mem[974] = 10'h1a4;
        mem[975] = 10'h28d;
        mem[976] = 10'h38b;
        mem[977] = 10'h213;
        mem[978] = 10'h23a;
        mem[979] = 10'h273;
        mem[980] = 10'h3b1;
        mem[981] = 10'h0c4;
        mem[982] = 10'h15b;
        mem[983] = 10'h057;
        mem[984] = 10'h0e2;
        mem[985] = 10'h1fe;
        mem[986] = 10'h22f;
        mem[987] = 10'h1db;
        mem[988] = 10'h248;
        mem[989] = 10'h36e;
        mem[990] = 10'h109;
        mem[991] = 10'h11e;
        mem[992] = 10'h2dc;
        mem[993] = 10'h265;
        mem[994] = 10'h34d;
        mem[995] = 10'h02b;
        mem[996] = 10'h111;
        mem[997] = 10'h37a;
        mem[998] = 10'h0c0;
        mem[999] = 10'h0ec;
        mem[1000] = 10'h341;
        mem[1001] = 10'h0f4;
        mem[1002] = 10'h088;
        mem[1003] = 10'h0cf;
        mem[1004] = 10'h237;
        mem[1005] = 10'h26a;
        mem[1006] = 10'h24f;
        mem[1007] = 10'h377;
        mem[1008] = 10'h35d;
        mem[1009] = 10'h1bf;
        mem[1010] = 10'h19b;
        mem[1011] = 10'h2bb;
        mem[1012] = 10'h0ff;
        mem[1013] = 10'h029;
        mem[1014] = 10'h247;
        mem[1015] = 10'h33d;
        mem[1016] = 10'h0f7;
        mem[1017] = 10'h383;
        mem[1018] = 10'h3ad;
        mem[1019] = 10'h1e3;
        mem[1020] = 10'h26d;
        mem[1021] = 10'h167;
        mem[1022] = 10'h1cd;
        mem[1023] = 10'h25f;
    end
endmodule

module odo_sbox_large6(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h185;
        mem[1] = 10'h2e3;
        mem[2] = 10'h352;
        mem[3] = 10'h04e;
        mem[4] = 10'h13f;
        mem[5] = 10'h3ab;
        mem[6] = 10'h1ac;
        mem[7] = 10'h04f;
        mem[8] = 10'h208;
        mem[9] = 10'h100;
        mem[10] = 10'h133;
        mem[11] = 10'h217;
        mem[12] = 10'h283;
        mem[13] = 10'h26f;
        mem[14] = 10'h380;
        mem[15] = 10'h1aa;
        mem[16] = 10'h12f;
        mem[17] = 10'h032;
        mem[18] = 10'h348;
        mem[19] = 10'h018;
        mem[20] = 10'h14a;
        mem[21] = 10'h00c;
        mem[22] = 10'h1a4;
        mem[23] = 10'h36a;
        mem[24] = 10'h039;
        mem[25] = 10'h2aa;
        mem[26] = 10'h0e2;
        mem[27] = 10'h04d;
        mem[28] = 10'h221;
        mem[29] = 10'h269;
        mem[30] = 10'h0f6;
        mem[31] = 10'h071;
        mem[32] = 10'h25a;
        mem[33] = 10'h08b;
        mem[34] = 10'h16a;
        mem[35] = 10'h37f;
        mem[36] = 10'h042;
        mem[37] = 10'h13b;
        mem[38] = 10'h132;
        mem[39] = 10'h122;
        mem[40] = 10'h026;
        mem[41] = 10'h059;
        mem[42] = 10'h3dd;
        mem[43] = 10'h1cb;
        mem[44] = 10'h070;
        mem[45] = 10'h3d1;
        mem[46] = 10'h229;
        mem[47] = 10'h3e6;
        mem[48] = 10'h0ea;
        mem[49] = 10'h3df;
        mem[50] = 10'h153;
        mem[51] = 10'h0b5;
        mem[52] = 10'h2da;
        mem[53] = 10'h0c1;
        mem[54] = 10'h11e;
        mem[55] = 10'h32f;
        mem[56] = 10'h0df;
        mem[57] = 10'h233;
        mem[58] = 10'h334;
        mem[59] = 10'h086;
        mem[60] = 10'h25c;
        mem[61] = 10'h073;
        mem[62] = 10'h2ce;
        mem[63] = 10'h004;
        mem[64] = 10'h06a;
        mem[65] = 10'h277;
        mem[66] = 10'h054;
        mem[67] = 10'h0b9;
        mem[68] = 10'h19c;
        mem[69] = 10'h1f9;
        mem[70] = 10'h323;
        mem[71] = 10'h0a5;
        mem[72] = 10'h16f;
        mem[73] = 10'h21d;
        mem[74] = 10'h24d;
        mem[75] = 10'h265;
        mem[76] = 10'h1f0;
        mem[77] = 10'h384;
        mem[78] = 10'h0f3;
        mem[79] = 10'h3db;
        mem[80] = 10'h0f4;
        mem[81] = 10'h25e;
        mem[82] = 10'h34c;
        mem[83] = 10'h046;
        mem[84] = 10'h0f8;
        mem[85] = 10'h0bf;
        mem[86] = 10'h168;
        mem[87] = 10'h095;
        mem[88] = 10'h3da;
        mem[89] = 10'h087;
        mem[90] = 10'h1d3;
        mem[91] = 10'h1fe;
        mem[92] = 10'h393;
        mem[93] = 10'h251;
        mem[94] = 10'h325;
        mem[95] = 10'h33a;
        mem[96] = 10'h276;
        mem[97] = 10'h302;
        mem[98] = 10'h023;
        mem[99] = 10'h2ca;
        mem[100] = 10'h1dd;
        mem[101] = 10'h3d0;
        mem[102] = 10'h117;
        mem[103] = 10'h19b;
        mem[104] = 10'h2f8;
        mem[105] = 10'h353;
        mem[106] = 10'h291;
        mem[107] = 10'h0cf;
        mem[108] = 10'h10f;
        mem[109] = 10'h306;
        mem[110] = 10'h374;
        mem[111] = 10'h088;
        mem[112] = 10'h252;
        mem[113] = 10'h18d;
        mem[114] = 10'h20d;
        mem[115] = 10'h224;
        mem[116] = 10'h378;
        mem[117] = 10'h21c;
        mem[118] = 10'h079;
        mem[119] = 10'h2dc;
        mem[120] = 10'h376;
        mem[121] = 10'h219;
        mem[122] = 10'h3e4;
        mem[123] = 10'h336;
        mem[124] = 10'h315;
        mem[125] = 10'h00e;
        mem[126] = 10'h0d5;
        mem[127] = 10'h395;
        mem[128] = 10'h199;
        mem[129] = 10'h0c2;
        mem[130] = 10'h1e6;
        mem[131] = 10'h2f5;
        mem[132] = 10'h090;
        mem[133] = 10'h1b0;
        mem[134] = 10'h07f;
        mem[135] = 10'h31e;
        mem[136] = 10'h15d;
        mem[137] = 10'h08d;
        mem[138] = 10'h1f4;
        mem[139] = 10'h147;
        mem[140] = 10'h170;
        mem[141] = 10'h181;
        mem[142] = 10'h1c3;
        mem[143] = 10'h267;
        mem[144] = 10'h0d7;
        mem[145] = 10'h2f2;
        mem[146] = 10'h189;
        mem[147] = 10'h379;
        mem[148] = 10'h17d;
        mem[149] = 10'h091;
        mem[150] = 10'h255;
        mem[151] = 10'h04c;
        mem[152] = 10'h161;
        mem[153] = 10'h27f;
        mem[154] = 10'h372;
        mem[155] = 10'h001;
        mem[156] = 10'h113;
        mem[157] = 10'h0b3;
        mem[158] = 10'h2e1;
        mem[159] = 10'h0bb;
        mem[160] = 10'h0ba;
        mem[161] = 10'h000;
        mem[162] = 10'h0d1;
        mem[163] = 10'h120;
        mem[164] = 10'h08f;
        mem[165] = 10'h207;
        mem[166] = 10'h078;
        mem[167] = 10'h0ac;
        mem[168] = 10'h3c1;
        mem[169] = 10'h10a;
        mem[170] = 10'h390;
        mem[171] = 10'h36b;
        mem[172] = 10'h005;
        mem[173] = 10'h3f3;
        mem[174] = 10'h3e5;
        mem[175] = 10'h215;
        mem[176] = 10'h32e;
        mem[177] = 10'h09d;
        mem[178] = 10'h263;
        mem[179] = 10'h1a6;
        mem[180] = 10'h33b;
        mem[181] = 10'h3c4;
        mem[182] = 10'h3ac;
        mem[183] = 10'h1b7;
        mem[184] = 10'h274;
        mem[185] = 10'h0c4;
        mem[186] = 10'h36e;
        mem[187] = 10'h313;
        mem[188] = 10'h21b;
        mem[189] = 10'h264;
        mem[190] = 10'h02c;
        mem[191] = 10'h3bf;
        mem[192] = 10'h1c6;
        mem[193] = 10'h114;
        mem[194] = 10'h15b;
        mem[195] = 10'h3c5;
        mem[196] = 10'h3ce;
        mem[197] = 10'h39f;
        mem[198] = 10'h301;
        mem[199] = 10'h3a6;
        mem[200] = 10'h103;
        mem[201] = 10'h319;
        mem[202] = 10'h27c;
        mem[203] = 10'h072;
        mem[204] = 10'h2db;
        mem[205] = 10'h0f7;
        mem[206] = 10'h3ad;
        mem[207] = 10'h0ec;
        mem[208] = 10'h1b4;
        mem[209] = 10'h36d;
        mem[210] = 10'h195;
        mem[211] = 10'h388;
        mem[212] = 10'h28f;
        mem[213] = 10'h055;
        mem[214] = 10'h299;
        mem[215] = 10'h06f;
        mem[216] = 10'h3ae;
        mem[217] = 10'h136;
        mem[218] = 10'h371;
        mem[219] = 10'h3f6;
        mem[220] = 10'h253;
        mem[221] = 10'h2c1;
        mem[222] = 10'h06b;
        mem[223] = 10'h068;
        mem[224] = 10'h2d8;
        mem[225] = 10'h3a3;
        mem[226] = 10'h037;
        mem[227] = 10'h3d6;
        mem[228] = 10'h31f;
        mem[229] = 10'h0ae;
        mem[230] = 10'h1f3;
        mem[231] = 10'h03d;
        mem[232] = 10'h2ae;
        mem[233] = 10'h02b;
        mem[234] = 10'h2fc;
        mem[235] = 10'h27e;
        mem[236] = 10'h10c;
        mem[237] = 10'h17b;
        mem[238] = 10'h2f1;
        mem[239] = 10'h089;
        mem[240] = 10'h09a;
        mem[241] = 10'h344;
        mem[242] = 10'h19f;
        mem[243] = 10'h1a2;
        mem[244] = 10'h0f1;
        mem[245] = 10'h027;
        mem[246] = 10'h21e;
        mem[247] = 10'h07b;
        mem[248] = 10'h0e0;
        mem[249] = 10'h1cc;
        mem[250] = 10'h1d2;
        mem[251] = 10'h118;
        mem[252] = 10'h0c7;
        mem[253] = 10'h320;
        mem[254] = 10'h230;
        mem[255] = 10'h3b3;
        mem[256] = 10'h38e;
        mem[257] = 10'h0fb;
        mem[258] = 10'h26c;
        mem[259] = 10'h0ed;
        mem[260] = 10'h30f;
        mem[261] = 10'h3a2;
        mem[262] = 10'h143;
        mem[263] = 10'h34b;
        mem[264] = 10'h318;
        mem[265] = 10'h2f6;
        mem[266] = 10'h2fe;
        mem[267] = 10'h2a0;
        mem[268] = 10'h3ef;
        mem[269] = 10'h36f;
        mem[270] = 10'h10e;
        mem[271] = 10'h0b2;
        mem[272] = 10'h0da;
        mem[273] = 10'h27b;
        mem[274] = 10'h28a;
        mem[275] = 10'h1ca;
        mem[276] = 10'h2bc;
        mem[277] = 10'h1af;
        mem[278] = 10'h11a;
        mem[279] = 10'h157;
        mem[280] = 10'h326;
        mem[281] = 10'h2d6;
        mem[282] = 10'h05b;
        mem[283] = 10'h37a;
        mem[284] = 10'h206;
        mem[285] = 10'h272;
        mem[286] = 10'h37c;
        mem[287] = 10'h048;
        mem[288] = 10'h28c;
        mem[289] = 10'h35f;
        mem[290] = 10'h332;
        mem[291] = 10'h196;
        mem[292] = 10'h1d7;
        mem[293] = 10'h27d;
        mem[294] = 10'h24f;
        mem[295] = 10'h385;
        mem[296] = 10'h37e;
        mem[297] = 10'h3ca;
        mem[298] = 10'h2c5;
        mem[299] = 10'h148;
        mem[300] = 10'h127;
        mem[301] = 10'h220;
        mem[302] = 10'h359;
        mem[303] = 10'h033;
        mem[304] = 10'h1eb;
        mem[305] = 10'h151;
        mem[306] = 10'h024;
        mem[307] = 10'h121;
        mem[308] = 10'h294;
        mem[309] = 10'h292;
        mem[310] = 10'h355;
        mem[311] = 10'h028;
        mem[312] = 10'h3fa;
        mem[313] = 10'h297;
        mem[314] = 10'h022;
        mem[315] = 10'h296;
        mem[316] = 10'h1f1;
        mem[317] = 10'h1fa;
        mem[318] = 10'h305;
        mem[319] = 10'h2de;
        mem[320] = 10'h099;
        mem[321] = 10'h00b;
        mem[322] = 10'h1d1;
        mem[323] = 10'h357;
        mem[324] = 10'h1bb;
        mem[325] = 10'h193;
        mem[326] = 10'h14e;
        mem[327] = 10'h1c2;
        mem[328] = 10'h2b7;
        mem[329] = 10'h210;
        mem[330] = 10'h084;
        mem[331] = 10'h2b3;
        mem[332] = 10'h298;
        mem[333] = 10'h07a;
        mem[334] = 10'h01d;
        mem[335] = 10'h3cf;
        mem[336] = 10'h1f7;
        mem[337] = 10'h04a;
        mem[338] = 10'h173;
        mem[339] = 10'h381;
        mem[340] = 10'h3f4;
        mem[341] = 10'h058;
        mem[342] = 10'h2e7;
        mem[343] = 10'h31b;
        mem[344] = 10'h234;
        mem[345] = 10'h14b;
        mem[346] = 10'h399;
        mem[347] = 10'h18e;
        mem[348] = 10'h149;
        mem[349] = 10'h0eb;
        mem[350] = 10'h1de;
        mem[351] = 10'h322;
        mem[352] = 10'h1a3;
        mem[353] = 10'h308;
        mem[354] = 10'h238;
        mem[355] = 10'h183;
        mem[356] = 10'h1e5;
        mem[357] = 10'h37b;
        mem[358] = 10'h050;
        mem[359] = 10'h281;
        mem[360] = 10'h202;
        mem[361] = 10'h0c0;
        mem[362] = 10'h130;
        mem[363] = 10'h32c;
        mem[364] = 10'h0aa;
        mem[365] = 10'h03e;
        mem[366] = 10'h16d;
        mem[367] = 10'h3a1;
        mem[368] = 10'h3fb;
        mem[369] = 10'h008;
        mem[370] = 10'h25f;
        mem[371] = 10'h0e6;
        mem[372] = 10'h1e2;
        mem[373] = 10'h167;
        mem[374] = 10'h2df;
        mem[375] = 10'h245;
        mem[376] = 10'h275;
        mem[377] = 10'h3f2;
        mem[378] = 10'h085;
        mem[379] = 10'h2e4;
        mem[380] = 10'h0f9;
        mem[381] = 10'h3c8;
        mem[382] = 10'h174;
        mem[383] = 10'h34a;
        mem[384] = 10'h16c;
        mem[385] = 10'h158;
        mem[386] = 10'h3bc;
        mem[387] = 10'h1db;
        mem[388] = 10'h11b;
        mem[389] = 10'h1d5;
        mem[390] = 10'h083;
        mem[391] = 10'h3f0;
        mem[392] = 10'h3be;
        mem[393] = 10'h007;
        mem[394] = 10'h18f;
        mem[395] = 10'h3b4;
        mem[396] = 10'h2e0;
        mem[397] = 10'h011;
        mem[398] = 10'h2fa;
        mem[399] = 10'h2b0;
        mem[400] = 10'h1c0;
        mem[401] = 10'h0cd;
        mem[402] = 10'h287;
        mem[403] = 10'h02a;
        mem[404] = 10'h2c8;
        mem[405] = 10'h080;
        mem[406] = 10'h159;
        mem[407] = 10'h171;
        mem[408] = 10'h2ad;
        mem[409] = 10'h389;
        mem[410] = 10'h289;
        mem[411] = 10'h10b;
        mem[412] = 10'h22b;
        mem[413] = 10'h06d;
        mem[414] = 10'h092;
        mem[415] = 10'h396;
        mem[416] = 10'h0cc;
        mem[417] = 10'h1c4;
        mem[418] = 10'h0b6;
        mem[419] = 10'h2af;
        mem[420] = 10'h284;
        mem[421] = 10'h2b8;
        mem[422] = 10'h12b;
        mem[423] = 10'h061;
        mem[424] = 10'h1a8;
        mem[425] = 10'h106;
        mem[426] = 10'h340;
        mem[427] = 10'h128;
        mem[428] = 10'h0c6;
        mem[429] = 10'h3af;
        mem[430] = 10'h31a;
        mem[431] = 10'h248;
        mem[432] = 10'h33e;
        mem[433] = 10'h107;
        mem[434] = 10'h1c5;
        mem[435] = 10'h0d8;
        mem[436] = 10'h1fd;
        mem[437] = 10'h386;
        mem[438] = 10'h1dc;
        mem[439] = 10'h0fd;
        mem[440] = 10'h329;
        mem[441] = 10'h169;
        mem[442] = 10'h134;
        mem[443] = 10'h0d4;
        mem[444] = 10'h2fd;
        mem[445] = 10'h250;
        mem[446] = 10'h266;
        mem[447] = 10'h34d;
        mem[448] = 10'h131;
        mem[449] = 10'h33c;
        mem[450] = 10'h2dd;
        mem[451] = 10'h017;
        mem[452] = 10'h278;
        mem[453] = 10'h119;
        mem[454] = 10'h01a;
        mem[455] = 10'h2eb;
        mem[456] = 10'h27a;
        mem[457] = 10'h21a;
        mem[458] = 10'h375;
        mem[459] = 10'h1b8;
        mem[460] = 10'h29c;
        mem[461] = 10'h0b1;
        mem[462] = 10'h163;
        mem[463] = 10'h066;
        mem[464] = 10'h2d3;
        mem[465] = 10'h38c;
        mem[466] = 10'h19d;
        mem[467] = 10'h249;
        mem[468] = 10'h162;
        mem[469] = 10'h1f5;
        mem[470] = 10'h3d7;
        mem[471] = 10'h057;
        mem[472] = 10'h1ae;
        mem[473] = 10'h043;
        mem[474] = 10'h38b;
        mem[475] = 10'h020;
        mem[476] = 10'h2ec;
        mem[477] = 10'h0fc;
        mem[478] = 10'h0af;
        mem[479] = 10'h138;
        mem[480] = 10'h0b0;
        mem[481] = 10'h26d;
        mem[482] = 10'h1b2;
        mem[483] = 10'h17c;
        mem[484] = 10'h0f2;
        mem[485] = 10'h09c;
        mem[486] = 10'h177;
        mem[487] = 10'h3fd;
        mem[488] = 10'h2bb;
        mem[489] = 10'h3bb;
        mem[490] = 10'h14f;
        mem[491] = 10'h341;
        mem[492] = 10'h0d2;
        mem[493] = 10'h13c;
        mem[494] = 10'h03b;
        mem[495] = 10'h17e;
        mem[496] = 10'h0b4;
        mem[497] = 10'h176;
        mem[498] = 10'h07d;
        mem[499] = 10'h2ac;
        mem[500] = 10'h20e;
        mem[501] = 10'h145;
        mem[502] = 10'h2d4;
        mem[503] = 10'h2fb;
        mem[504] = 10'h223;
        mem[505] = 10'h097;
        mem[506] = 10'h2b5;
        mem[507] = 10'h1d4;
        mem[508] = 10'h349;
        mem[509] = 10'h21f;
        mem[510] = 10'h293;
        mem[511] = 10'h38d;
        mem[512] = 10'h373;
        mem[513] = 10'h3d3;
        mem[514] = 10'h3fe;
        mem[515] = 10'h3de;
        mem[516] = 10'h09e;
        mem[517] = 10'h240;
        mem[518] = 10'h342;
        mem[519] = 10'h2cd;
        mem[520] = 10'h182;
        mem[521] = 10'h261;
        mem[522] = 10'h262;
        mem[523] = 10'h104;
        mem[524] = 10'h2ee;
        mem[525] = 10'h0ff;
        mem[526] = 10'h1f6;
        mem[527] = 10'h08a;
        mem[528] = 10'h34f;
        mem[529] = 10'h377;
        mem[530] = 10'h232;
        mem[531] = 10'h20b;
        mem[532] = 10'h04b;
        mem[533] = 10'h0ce;
        mem[534] = 10'h05c;
        mem[535] = 10'h26b;
        mem[536] = 10'h257;
        mem[537] = 10'h0fa;
        mem[538] = 10'h3e8;
        mem[539] = 10'h346;
        mem[540] = 10'h082;
        mem[541] = 10'h1e3;
        mem[542] = 10'h175;
        mem[543] = 10'h350;
        mem[544] = 10'h08e;
        mem[545] = 10'h309;
        mem[546] = 10'h015;
        mem[547] = 10'h200;
        mem[548] = 10'h3fc;
        mem[549] = 10'h2c0;
        mem[550] = 10'h1f2;
        mem[551] = 10'h338;
        mem[552] = 10'h035;
        mem[553] = 10'h178;
        mem[554] = 10'h144;
        mem[555] = 10'h35e;
        mem[556] = 10'h110;
        mem[557] = 10'h17a;
        mem[558] = 10'h18a;
        mem[559] = 10'h19a;
        mem[560] = 10'h156;
        mem[561] = 10'h002;
        mem[562] = 10'h2be;
        mem[563] = 10'h0a4;
        mem[564] = 10'h0a8;
        mem[565] = 10'h146;
        mem[566] = 10'h3ed;
        mem[567] = 10'h12d;
        mem[568] = 10'h139;
        mem[569] = 10'h019;
        mem[570] = 10'h0e5;
        mem[571] = 10'h26a;
        mem[572] = 10'h062;
        mem[573] = 10'h135;
        mem[574] = 10'h1ec;
        mem[575] = 10'h28d;
        mem[576] = 10'h3a5;
        mem[577] = 10'h129;
        mem[578] = 10'h188;
        mem[579] = 10'h2f4;
        mem[580] = 10'h2ba;
        mem[581] = 10'h31c;
        mem[582] = 10'h3b9;
        mem[583] = 10'h094;
        mem[584] = 10'h105;
        mem[585] = 10'h13e;
        mem[586] = 10'h23c;
        mem[587] = 10'h1c9;
        mem[588] = 10'h10d;
        mem[589] = 10'h239;
        mem[590] = 10'h3f5;
        mem[591] = 10'h112;
        mem[592] = 10'h1c7;
        mem[593] = 10'h1e1;
        mem[594] = 10'h369;
        mem[595] = 10'h0a6;
        mem[596] = 10'h0e7;
        mem[597] = 10'h2cb;
        mem[598] = 10'h09b;
        mem[599] = 10'h3a0;
        mem[600] = 10'h23a;
        mem[601] = 10'h337;
        mem[602] = 10'h02f;
        mem[603] = 10'h3b8;
        mem[604] = 10'h165;
        mem[605] = 10'h339;
        mem[606] = 10'h30a;
        mem[607] = 10'h211;
        mem[608] = 10'h140;
        mem[609] = 10'h22a;
        mem[610] = 10'h0d6;
        mem[611] = 10'h394;
        mem[612] = 10'h0d0;
        mem[613] = 10'h3ee;
        mem[614] = 10'h398;
        mem[615] = 10'h222;
        mem[616] = 10'h35b;
        mem[617] = 10'h180;
        mem[618] = 10'h24b;
        mem[619] = 10'h152;
        mem[620] = 10'h29e;
        mem[621] = 10'h172;
        mem[622] = 10'h333;
        mem[623] = 10'h2c4;
        mem[624] = 10'h2f7;
        mem[625] = 10'h14d;
        mem[626] = 10'h191;
        mem[627] = 10'h331;
        mem[628] = 10'h345;
        mem[629] = 10'h101;
        mem[630] = 10'h081;
        mem[631] = 10'h2e6;
        mem[632] = 10'h2b1;
        mem[633] = 10'h204;
        mem[634] = 10'h242;
        mem[635] = 10'h0a9;
        mem[636] = 10'h38a;
        mem[637] = 10'h01c;
        mem[638] = 10'h2e5;
        mem[639] = 10'h1e8;
        mem[640] = 10'h00a;
        mem[641] = 10'h2f9;
        mem[642] = 10'h2bd;
        mem[643] = 10'h247;
        mem[644] = 10'h360;
        mem[645] = 10'h150;
        mem[646] = 10'h15e;
        mem[647] = 10'h3d9;
        mem[648] = 10'h32b;
        mem[649] = 10'h307;
        mem[650] = 10'h286;
        mem[651] = 10'h370;
        mem[652] = 10'h2c3;
        mem[653] = 10'h198;
        mem[654] = 10'h347;
        mem[655] = 10'h2f3;
        mem[656] = 10'h216;
        mem[657] = 10'h164;
        mem[658] = 10'h051;
        mem[659] = 10'h227;
        mem[660] = 10'h0d9;
        mem[661] = 10'h351;
        mem[662] = 10'h01e;
        mem[663] = 10'h013;
        mem[664] = 10'h303;
        mem[665] = 10'h13a;
        mem[666] = 10'h2c2;
        mem[667] = 10'h154;
        mem[668] = 10'h2a3;
        mem[669] = 10'h0c9;
        mem[670] = 10'h3d4;
        mem[671] = 10'h064;
        mem[672] = 10'h0f0;
        mem[673] = 10'h056;
        mem[674] = 10'h3a9;
        mem[675] = 10'h07c;
        mem[676] = 10'h35c;
        mem[677] = 10'h01f;
        mem[678] = 10'h197;
        mem[679] = 10'h155;
        mem[680] = 10'h15c;
        mem[681] = 10'h271;
        mem[682] = 10'h1f8;
        mem[683] = 10'h08c;
        mem[684] = 10'h029;
        mem[685] = 10'h3ec;
        mem[686] = 10'h32d;
        mem[687] = 10'h3eb;
        mem[688] = 10'h016;
        mem[689] = 10'h214;
        mem[690] = 10'h1e0;
        mem[691] = 10'h368;
        mem[692] = 10'h39c;
        mem[693] = 10'h1e7;
        mem[694] = 10'h30b;
        mem[695] = 10'h225;
        mem[696] = 10'h1d8;
        mem[697] = 10'h0cb;
        mem[698] = 10'h3b5;
        mem[699] = 10'h096;
        mem[700] = 10'h021;
        mem[701] = 10'h22e;
        mem[702] = 10'h3dc;
        mem[703] = 10'h00f;
        mem[704] = 10'h14c;
        mem[705] = 10'h125;
        mem[706] = 10'h3cc;
        mem[707] = 10'h38f;
        mem[708] = 10'h2c9;
        mem[709] = 10'h282;
        mem[710] = 10'h0b7;
        mem[711] = 10'h12e;
        mem[712] = 10'h366;
        mem[713] = 10'h0a3;
        mem[714] = 10'h1ee;
        mem[715] = 10'h3b7;
        mem[716] = 10'h1ba;
        mem[717] = 10'h2d1;
        mem[718] = 10'h290;
        mem[719] = 10'h109;
        mem[720] = 10'h258;
        mem[721] = 10'h3c0;
        mem[722] = 10'h304;
        mem[723] = 10'h3f8;
        mem[724] = 10'h1d6;
        mem[725] = 10'h270;
        mem[726] = 10'h231;
        mem[727] = 10'h115;
        mem[728] = 10'h0a1;
        mem[729] = 10'h25b;
        mem[730] = 10'h142;
        mem[731] = 10'h382;
        mem[732] = 10'h365;
        mem[733] = 10'h1fc;
        mem[734] = 10'h383;
        mem[735] = 10'h2ff;
        mem[736] = 10'h02d;
        mem[737] = 10'h19e;
        mem[738] = 10'h012;
        mem[739] = 10'h1a0;
        mem[740] = 10'h237;
        mem[741] = 10'h22f;
        mem[742] = 10'h3cd;
        mem[743] = 10'h22d;
        mem[744] = 10'h0ef;
        mem[745] = 10'h2b4;
        mem[746] = 10'h23e;
        mem[747] = 10'h39a;
        mem[748] = 10'h3aa;
        mem[749] = 10'h025;
        mem[750] = 10'h15f;
        mem[751] = 10'h3e3;
        mem[752] = 10'h362;
        mem[753] = 10'h160;
        mem[754] = 10'h0ab;
        mem[755] = 10'h111;
        mem[756] = 10'h3c3;
        mem[757] = 10'h213;
        mem[758] = 10'h194;
        mem[759] = 10'h045;
        mem[760] = 10'h23d;
        mem[761] = 10'h367;
        mem[762] = 10'h2b9;
        mem[763] = 10'h328;
        mem[764] = 10'h030;
        mem[765] = 10'h0e4;
        mem[766] = 10'h218;
        mem[767] = 10'h23f;
        mem[768] = 10'h16e;
        mem[769] = 10'h321;
        mem[770] = 10'h074;
        mem[771] = 10'h39e;
        mem[772] = 10'h2d0;
        mem[773] = 10'h241;
        mem[774] = 10'h0dd;
        mem[775] = 10'h2ea;
        mem[776] = 10'h256;
        mem[777] = 10'h30c;
        mem[778] = 10'h00d;
        mem[779] = 10'h2e2;
        mem[780] = 10'h1bc;
        mem[781] = 10'h3f1;
        mem[782] = 10'h3f7;
        mem[783] = 10'h2ef;
        mem[784] = 10'h288;
        mem[785] = 10'h39d;
        mem[786] = 10'h1a9;
        mem[787] = 10'h39b;
        mem[788] = 10'h1d0;
        mem[789] = 10'h3a7;
        mem[790] = 10'h268;
        mem[791] = 10'h28e;
        mem[792] = 10'h0c3;
        mem[793] = 10'h392;
        mem[794] = 10'h327;
        mem[795] = 10'h041;
        mem[796] = 10'h391;
        mem[797] = 10'h1b1;
        mem[798] = 10'h2a6;
        mem[799] = 10'h3e0;
        mem[800] = 10'h01b;
        mem[801] = 10'h18c;
        mem[802] = 10'h1fb;
        mem[803] = 10'h0e8;
        mem[804] = 10'h358;
        mem[805] = 10'h05f;
        mem[806] = 10'h28b;
        mem[807] = 10'h098;
        mem[808] = 10'h31d;
        mem[809] = 10'h36c;
        mem[810] = 10'h24a;
        mem[811] = 10'h2a4;
        mem[812] = 10'h0bc;
        mem[813] = 10'h228;
        mem[814] = 10'h1b6;
        mem[815] = 10'h201;
        mem[816] = 10'h186;
        mem[817] = 10'h1ea;
        mem[818] = 10'h35d;
        mem[819] = 10'h141;
        mem[820] = 10'h209;
        mem[821] = 10'h1df;
        mem[822] = 10'h12c;
        mem[823] = 10'h2b2;
        mem[824] = 10'h02e;
        mem[825] = 10'h014;
        mem[826] = 10'h11d;
        mem[827] = 10'h3ea;
        mem[828] = 10'h2b6;
        mem[829] = 10'h2c7;
        mem[830] = 10'h1d9;
        mem[831] = 10'h3a4;
        mem[832] = 10'h361;
        mem[833] = 10'h184;
        mem[834] = 10'h12a;
        mem[835] = 10'h363;
        mem[836] = 10'h0de;
        mem[837] = 10'h37d;
        mem[838] = 10'h063;
        mem[839] = 10'h316;
        mem[840] = 10'h330;
        mem[841] = 10'h26e;
        mem[842] = 10'h3c7;
        mem[843] = 10'h006;
        mem[844] = 10'h1ce;
        mem[845] = 10'h1cd;
        mem[846] = 10'h010;
        mem[847] = 10'h0a7;
        mem[848] = 10'h05e;
        mem[849] = 10'h205;
        mem[850] = 10'h179;
        mem[851] = 10'h003;
        mem[852] = 10'h23b;
        mem[853] = 10'h047;
        mem[854] = 10'h285;
        mem[855] = 10'h11f;
        mem[856] = 10'h3ba;
        mem[857] = 10'h3d5;
        mem[858] = 10'h0ad;
        mem[859] = 10'h044;
        mem[860] = 10'h2a5;
        mem[861] = 10'h3b0;
        mem[862] = 10'h1bf;
        mem[863] = 10'h1e9;
        mem[864] = 10'h065;
        mem[865] = 10'h203;
        mem[866] = 10'h137;
        mem[867] = 10'h0a0;
        mem[868] = 10'h3d8;
        mem[869] = 10'h3cb;
        mem[870] = 10'h273;
        mem[871] = 10'h05d;
        mem[872] = 10'h3b2;
        mem[873] = 10'h077;
        mem[874] = 10'h335;
        mem[875] = 10'h246;
        mem[876] = 10'h311;
        mem[877] = 10'h1be;
        mem[878] = 10'h108;
        mem[879] = 10'h13d;
        mem[880] = 10'h1cf;
        mem[881] = 10'h038;
        mem[882] = 10'h2a8;
        mem[883] = 10'h2e8;
        mem[884] = 10'h11c;
        mem[885] = 10'h0ca;
        mem[886] = 10'h07e;
        mem[887] = 10'h300;
        mem[888] = 10'h33f;
        mem[889] = 10'h192;
        mem[890] = 10'h0e9;
        mem[891] = 10'h2c6;
        mem[892] = 10'h2a2;
        mem[893] = 10'h30e;
        mem[894] = 10'h310;
        mem[895] = 10'h3e2;
        mem[896] = 10'h0db;
        mem[897] = 10'h126;
        mem[898] = 10'h343;
        mem[899] = 10'h1a5;
        mem[900] = 10'h279;
        mem[901] = 10'h29b;
        mem[902] = 10'h067;
        mem[903] = 10'h2d9;
        mem[904] = 10'h226;
        mem[905] = 10'h009;
        mem[906] = 10'h16b;
        mem[907] = 10'h24e;
        mem[908] = 10'h397;
        mem[909] = 10'h2ed;
        mem[910] = 10'h387;
        mem[911] = 10'h354;
        mem[912] = 10'h3e9;
        mem[913] = 10'h29d;
        mem[914] = 10'h3c6;
        mem[915] = 10'h2d2;
        mem[916] = 10'h243;
        mem[917] = 10'h036;
        mem[918] = 10'h1ab;
        mem[919] = 10'h0c8;
        mem[920] = 10'h076;
        mem[921] = 10'h1a1;
        mem[922] = 10'h1da;
        mem[923] = 10'h18b;
        mem[924] = 10'h0b8;
        mem[925] = 10'h124;
        mem[926] = 10'h2a9;
        mem[927] = 10'h2cf;
        mem[928] = 10'h1b5;
        mem[929] = 10'h1a7;
        mem[930] = 10'h17f;
        mem[931] = 10'h3ff;
        mem[932] = 10'h093;
        mem[933] = 10'h034;
        mem[934] = 10'h0f5;
        mem[935] = 10'h259;
        mem[936] = 10'h03c;
        mem[937] = 10'h33d;
        mem[938] = 10'h3a8;
        mem[939] = 10'h3bd;
        mem[940] = 10'h30d;
        mem[941] = 10'h1c1;
        mem[942] = 10'h34e;
        mem[943] = 10'h3c9;
        mem[944] = 10'h35a;
        mem[945] = 10'h212;
        mem[946] = 10'h049;
        mem[947] = 10'h187;
        mem[948] = 10'h2cc;
        mem[949] = 10'h2d5;
        mem[950] = 10'h0a2;
        mem[951] = 10'h052;
        mem[952] = 10'h3f9;
        mem[953] = 10'h1ef;
        mem[954] = 10'h0ee;
        mem[955] = 10'h314;
        mem[956] = 10'h0c5;
        mem[957] = 10'h0d3;
        mem[958] = 10'h260;
        mem[959] = 10'h166;
        mem[960] = 10'h1ff;
        mem[961] = 10'h312;
        mem[962] = 10'h0bd;
        mem[963] = 10'h2f0;
        mem[964] = 10'h102;
        mem[965] = 10'h0be;
        mem[966] = 10'h3b6;
        mem[967] = 10'h05a;
        mem[968] = 10'h236;
        mem[969] = 10'h03f;
        mem[970] = 10'h06e;
        mem[971] = 10'h1ad;
        mem[972] = 10'h15a;
        mem[973] = 10'h244;
        mem[974] = 10'h0fe;
        mem[975] = 10'h116;
        mem[976] = 10'h29f;
        mem[977] = 10'h1bd;
        mem[978] = 10'h1b9;
        mem[979] = 10'h280;
        mem[980] = 10'h190;
        mem[981] = 10'h25d;
        mem[982] = 10'h0e3;
        mem[983] = 10'h24c;
        mem[984] = 10'h075;
        mem[985] = 10'h031;
        mem[986] = 10'h0e1;
        mem[987] = 10'h1c8;
        mem[988] = 10'h0dc;
        mem[989] = 10'h2e9;
        mem[990] = 10'h20a;
        mem[991] = 10'h32a;
        mem[992] = 10'h295;
        mem[993] = 10'h1ed;
        mem[994] = 10'h040;
        mem[995] = 10'h2bf;
        mem[996] = 10'h2a7;
        mem[997] = 10'h2d7;
        mem[998] = 10'h3d2;
        mem[999] = 10'h317;
        mem[1000] = 10'h356;
        mem[1001] = 10'h29a;
        mem[1002] = 10'h060;
        mem[1003] = 10'h235;
        mem[1004] = 10'h3e1;
        mem[1005] = 10'h364;
        mem[1006] = 10'h22c;
        mem[1007] = 10'h3b1;
        mem[1008] = 10'h324;
        mem[1009] = 10'h20f;
        mem[1010] = 10'h2a1;
        mem[1011] = 10'h03a;
        mem[1012] = 10'h3c2;
        mem[1013] = 10'h123;
        mem[1014] = 10'h069;
        mem[1015] = 10'h3e7;
        mem[1016] = 10'h20c;
        mem[1017] = 10'h2ab;
        mem[1018] = 10'h053;
        mem[1019] = 10'h254;
        mem[1020] = 10'h09f;
        mem[1021] = 10'h1b3;
        mem[1022] = 10'h1e4;
        mem[1023] = 10'h06c;
    end
endmodule

module odo_sbox_large7(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h112;
        mem[1] = 10'h2b2;
        mem[2] = 10'h04b;
        mem[3] = 10'h1b1;
        mem[4] = 10'h3c0;
        mem[5] = 10'h1e5;
        mem[6] = 10'h171;
        mem[7] = 10'h22c;
        mem[8] = 10'h10d;
        mem[9] = 10'h033;
        mem[10] = 10'h21e;
        mem[11] = 10'h08b;
        mem[12] = 10'h265;
        mem[13] = 10'h20f;
        mem[14] = 10'h2dc;
        mem[15] = 10'h147;
        mem[16] = 10'h2a1;
        mem[17] = 10'h064;
        mem[18] = 10'h33a;
        mem[19] = 10'h07f;
        mem[20] = 10'h1cc;
        mem[21] = 10'h19f;
        mem[22] = 10'h047;
        mem[23] = 10'h13b;
        mem[24] = 10'h1d5;
        mem[25] = 10'h1c4;
        mem[26] = 10'h004;
        mem[27] = 10'h27e;
        mem[28] = 10'h36e;
        mem[29] = 10'h246;
        mem[30] = 10'h09e;
        mem[31] = 10'h3d4;
        mem[32] = 10'h002;
        mem[33] = 10'h204;
        mem[34] = 10'h36c;
        mem[35] = 10'h0aa;
        mem[36] = 10'h270;
        mem[37] = 10'h341;
        mem[38] = 10'h035;
        mem[39] = 10'h345;
        mem[40] = 10'h250;
        mem[41] = 10'h322;
        mem[42] = 10'h049;
        mem[43] = 10'h3e6;
        mem[44] = 10'h24c;
        mem[45] = 10'h173;
        mem[46] = 10'h29a;
        mem[47] = 10'h244;
        mem[48] = 10'h0fd;
        mem[49] = 10'h3fe;
        mem[50] = 10'h15b;
        mem[51] = 10'h229;
        mem[52] = 10'h242;
        mem[53] = 10'h1c0;
        mem[54] = 10'h261;
        mem[55] = 10'h351;
        mem[56] = 10'h383;
        mem[57] = 10'h02d;
        mem[58] = 10'h2ea;
        mem[59] = 10'h190;
        mem[60] = 10'h099;
        mem[61] = 10'h0b1;
        mem[62] = 10'h25f;
        mem[63] = 10'h2c9;
        mem[64] = 10'h3fd;
        mem[65] = 10'h2f9;
        mem[66] = 10'h249;
        mem[67] = 10'h368;
        mem[68] = 10'h135;
        mem[69] = 10'h018;
        mem[70] = 10'h32b;
        mem[71] = 10'h104;
        mem[72] = 10'h014;
        mem[73] = 10'h199;
        mem[74] = 10'h037;
        mem[75] = 10'h36b;
        mem[76] = 10'h366;
        mem[77] = 10'h146;
        mem[78] = 10'h20e;
        mem[79] = 10'h3d2;
        mem[80] = 10'h303;
        mem[81] = 10'h3c5;
        mem[82] = 10'h1af;
        mem[83] = 10'h2ee;
        mem[84] = 10'h3e3;
        mem[85] = 10'h3f3;
        mem[86] = 10'h081;
        mem[87] = 10'h178;
        mem[88] = 10'h073;
        mem[89] = 10'h0d8;
        mem[90] = 10'h048;
        mem[91] = 10'h34d;
        mem[92] = 10'h2b8;
        mem[93] = 10'h293;
        mem[94] = 10'h34f;
        mem[95] = 10'h3da;
        mem[96] = 10'h35a;
        mem[97] = 10'h0e1;
        mem[98] = 10'h1fd;
        mem[99] = 10'h332;
        mem[100] = 10'h077;
        mem[101] = 10'h23a;
        mem[102] = 10'h335;
        mem[103] = 10'h355;
        mem[104] = 10'h16e;
        mem[105] = 10'h16f;
        mem[106] = 10'h3ca;
        mem[107] = 10'h3c7;
        mem[108] = 10'h352;
        mem[109] = 10'h105;
        mem[110] = 10'h0f6;
        mem[111] = 10'h2ef;
        mem[112] = 10'h096;
        mem[113] = 10'h0e5;
        mem[114] = 10'h35e;
        mem[115] = 10'h0dd;
        mem[116] = 10'h21c;
        mem[117] = 10'h0e6;
        mem[118] = 10'h307;
        mem[119] = 10'h1c9;
        mem[120] = 10'h2a2;
        mem[121] = 10'h084;
        mem[122] = 10'h31e;
        mem[123] = 10'h039;
        mem[124] = 10'h310;
        mem[125] = 10'h1d4;
        mem[126] = 10'h211;
        mem[127] = 10'h2a0;
        mem[128] = 10'h272;
        mem[129] = 10'h0f1;
        mem[130] = 10'h11b;
        mem[131] = 10'h1bc;
        mem[132] = 10'h0ac;
        mem[133] = 10'h0e7;
        mem[134] = 10'h155;
        mem[135] = 10'h143;
        mem[136] = 10'h33f;
        mem[137] = 10'h0ce;
        mem[138] = 10'h362;
        mem[139] = 10'h208;
        mem[140] = 10'h0f5;
        mem[141] = 10'h03f;
        mem[142] = 10'h1e1;
        mem[143] = 10'h1b7;
        mem[144] = 10'h0d3;
        mem[145] = 10'h311;
        mem[146] = 10'h2b7;
        mem[147] = 10'h06e;
        mem[148] = 10'h393;
        mem[149] = 10'h39c;
        mem[150] = 10'h3be;
        mem[151] = 10'h226;
        mem[152] = 10'h21b;
        mem[153] = 10'h060;
        mem[154] = 10'h1b6;
        mem[155] = 10'h168;
        mem[156] = 10'h00a;
        mem[157] = 10'h3a9;
        mem[158] = 10'h34e;
        mem[159] = 10'h03b;
        mem[160] = 10'h215;
        mem[161] = 10'h15a;
        mem[162] = 10'h140;
        mem[163] = 10'h3f1;
        mem[164] = 10'h2c1;
        mem[165] = 10'h327;
        mem[166] = 10'h006;
        mem[167] = 10'h0cc;
        mem[168] = 10'h31d;
        mem[169] = 10'h13c;
        mem[170] = 10'h016;
        mem[171] = 10'h259;
        mem[172] = 10'h2f2;
        mem[173] = 10'h283;
        mem[174] = 10'h0c6;
        mem[175] = 10'h2d6;
        mem[176] = 10'h3b2;
        mem[177] = 10'h2fe;
        mem[178] = 10'h052;
        mem[179] = 10'h37e;
        mem[180] = 10'h24b;
        mem[181] = 10'h1de;
        mem[182] = 10'h1c7;
        mem[183] = 10'h3c3;
        mem[184] = 10'h1ae;
        mem[185] = 10'h34a;
        mem[186] = 10'h0ff;
        mem[187] = 10'h2d9;
        mem[188] = 10'h262;
        mem[189] = 10'h18a;
        mem[190] = 10'h336;
        mem[191] = 10'h0fb;
        mem[192] = 10'h225;
        mem[193] = 10'h041;
        mem[194] = 10'h16a;
        mem[195] = 10'h2e3;
        mem[196] = 10'h378;
        mem[197] = 10'h3c9;
        mem[198] = 10'h11a;
        mem[199] = 10'h0c1;
        mem[200] = 10'h3f0;
        mem[201] = 10'h0e4;
        mem[202] = 10'h278;
        mem[203] = 10'h297;
        mem[204] = 10'h062;
        mem[205] = 10'h0c4;
        mem[206] = 10'h18e;
        mem[207] = 10'h36a;
        mem[208] = 10'h0a1;
        mem[209] = 10'h299;
        mem[210] = 10'h19e;
        mem[211] = 10'h069;
        mem[212] = 10'h2f8;
        mem[213] = 10'h032;
        mem[214] = 10'h31c;
        mem[215] = 10'h291;
        mem[216] = 10'h23c;
        mem[217] = 10'h388;
        mem[218] = 10'h1b8;
        mem[219] = 10'h083;
        mem[220] = 10'h09b;
        mem[221] = 10'h2fc;
        mem[222] = 10'h119;
        mem[223] = 10'h3fc;
        mem[224] = 10'h2be;
        mem[225] = 10'h114;
        mem[226] = 10'h397;
        mem[227] = 10'h38d;
        mem[228] = 10'h3e7;
        mem[229] = 10'h093;
        mem[230] = 10'h0a8;
        mem[231] = 10'h28e;
        mem[232] = 10'h0bc;
        mem[233] = 10'h2cc;
        mem[234] = 10'h3db;
        mem[235] = 10'h139;
        mem[236] = 10'h254;
        mem[237] = 10'h13f;
        mem[238] = 10'h36f;
        mem[239] = 10'h370;
        mem[240] = 10'h124;
        mem[241] = 10'h217;
        mem[242] = 10'h0de;
        mem[243] = 10'h053;
        mem[244] = 10'h1f9;
        mem[245] = 10'h380;
        mem[246] = 10'h136;
        mem[247] = 10'h201;
        mem[248] = 10'h315;
        mem[249] = 10'h28c;
        mem[250] = 10'h2d4;
        mem[251] = 10'h19b;
        mem[252] = 10'h38f;
        mem[253] = 10'h076;
        mem[254] = 10'h24d;
        mem[255] = 10'h1e8;
        mem[256] = 10'h2f3;
        mem[257] = 10'h3f9;
        mem[258] = 10'h26d;
        mem[259] = 10'h32c;
        mem[260] = 10'h15d;
        mem[261] = 10'h2c7;
        mem[262] = 10'h2bc;
        mem[263] = 10'h10f;
        mem[264] = 10'h0d6;
        mem[265] = 10'h3f5;
        mem[266] = 10'h288;
        mem[267] = 10'h090;
        mem[268] = 10'h05e;
        mem[269] = 10'h1ec;
        mem[270] = 10'h07c;
        mem[271] = 10'h0be;
        mem[272] = 10'h234;
        mem[273] = 10'h138;
        mem[274] = 10'h141;
        mem[275] = 10'h2d8;
        mem[276] = 10'h3f4;
        mem[277] = 10'h240;
        mem[278] = 10'h0ef;
        mem[279] = 10'h1d7;
        mem[280] = 10'h188;
        mem[281] = 10'h309;
        mem[282] = 10'h3dc;
        mem[283] = 10'h2c8;
        mem[284] = 10'h275;
        mem[285] = 10'h106;
        mem[286] = 10'h339;
        mem[287] = 10'h1a2;
        mem[288] = 10'h06b;
        mem[289] = 10'h120;
        mem[290] = 10'h1b4;
        mem[291] = 10'h359;
        mem[292] = 10'h364;
        mem[293] = 10'h245;
        mem[294] = 10'h198;
        mem[295] = 10'h255;
        mem[296] = 10'h1f1;
        mem[297] = 10'h2ca;
        mem[298] = 10'h2c2;
        mem[299] = 10'h323;
        mem[300] = 10'h03d;
        mem[301] = 10'h213;
        mem[302] = 10'h103;
        mem[303] = 10'h239;
        mem[304] = 10'h28a;
        mem[305] = 10'h02f;
        mem[306] = 10'h3a6;
        mem[307] = 10'h2f4;
        mem[308] = 10'h02e;
        mem[309] = 10'h286;
        mem[310] = 10'h3f6;
        mem[311] = 10'h264;
        mem[312] = 10'h27b;
        mem[313] = 10'h251;
        mem[314] = 10'h333;
        mem[315] = 10'h019;
        mem[316] = 10'h2e4;
        mem[317] = 10'h3d1;
        mem[318] = 10'h266;
        mem[319] = 10'h1fa;
        mem[320] = 10'h306;
        mem[321] = 10'h330;
        mem[322] = 10'h04d;
        mem[323] = 10'h2b1;
        mem[324] = 10'h2bf;
        mem[325] = 10'h063;
        mem[326] = 10'h14a;
        mem[327] = 10'h0d2;
        mem[328] = 10'h2f1;
        mem[329] = 10'h0e9;
        mem[330] = 10'h361;
        mem[331] = 10'h2da;
        mem[332] = 10'h1db;
        mem[333] = 10'h2cf;
        mem[334] = 10'h06c;
        mem[335] = 10'h3a5;
        mem[336] = 10'h27a;
        mem[337] = 10'h30e;
        mem[338] = 10'h3d7;
        mem[339] = 10'h21a;
        mem[340] = 10'h100;
        mem[341] = 10'h3b3;
        mem[342] = 10'h36d;
        mem[343] = 10'h209;
        mem[344] = 10'h0ea;
        mem[345] = 10'h39a;
        mem[346] = 10'h1ad;
        mem[347] = 10'h3cc;
        mem[348] = 10'h3e8;
        mem[349] = 10'h13e;
        mem[350] = 10'h38c;
        mem[351] = 10'h373;
        mem[352] = 10'h17d;
        mem[353] = 10'h12d;
        mem[354] = 10'h20a;
        mem[355] = 10'h0a2;
        mem[356] = 10'h01b;
        mem[357] = 10'h1ce;
        mem[358] = 10'h1f8;
        mem[359] = 10'h06f;
        mem[360] = 10'h102;
        mem[361] = 10'h25d;
        mem[362] = 10'h03a;
        mem[363] = 10'h2d0;
        mem[364] = 10'h329;
        mem[365] = 10'h023;
        mem[366] = 10'h055;
        mem[367] = 10'h03e;
        mem[368] = 10'h30d;
        mem[369] = 10'h017;
        mem[370] = 10'h256;
        mem[371] = 10'h31b;
        mem[372] = 10'h034;
        mem[373] = 10'h2b5;
        mem[374] = 10'h237;
        mem[375] = 10'h221;
        mem[376] = 10'h0ca;
        mem[377] = 10'h010;
        mem[378] = 10'h061;
        mem[379] = 10'h13a;
        mem[380] = 10'h07e;
        mem[381] = 10'h074;
        mem[382] = 10'h013;
        mem[383] = 10'h3d5;
        mem[384] = 10'h26c;
        mem[385] = 10'h194;
        mem[386] = 10'h3d0;
        mem[387] = 10'h14e;
        mem[388] = 10'h11e;
        mem[389] = 10'h00d;
        mem[390] = 10'h0a3;
        mem[391] = 10'h027;
        mem[392] = 10'h2c6;
        mem[393] = 10'h046;
        mem[394] = 10'h319;
        mem[395] = 10'h282;
        mem[396] = 10'h17f;
        mem[397] = 10'h117;
        mem[398] = 10'h2b6;
        mem[399] = 10'h285;
        mem[400] = 10'h223;
        mem[401] = 10'h38b;
        mem[402] = 10'h091;
        mem[403] = 10'h34c;
        mem[404] = 10'h3de;
        mem[405] = 10'h0b4;
        mem[406] = 10'h17b;
        mem[407] = 10'h180;
        mem[408] = 10'h15c;
        mem[409] = 10'h142;
        mem[410] = 10'h3ba;
        mem[411] = 10'h353;
        mem[412] = 10'h3c2;
        mem[413] = 10'h07d;
        mem[414] = 10'h3fb;
        mem[415] = 10'h268;
        mem[416] = 10'h044;
        mem[417] = 10'h321;
        mem[418] = 10'h342;
        mem[419] = 10'h236;
        mem[420] = 10'h3a8;
        mem[421] = 10'h23d;
        mem[422] = 10'h358;
        mem[423] = 10'h2a9;
        mem[424] = 10'h3cd;
        mem[425] = 10'h350;
        mem[426] = 10'h01c;
        mem[427] = 10'h0c2;
        mem[428] = 10'h273;
        mem[429] = 10'h0f2;
        mem[430] = 10'h2c3;
        mem[431] = 10'h148;
        mem[432] = 10'h2e7;
        mem[433] = 10'h33e;
        mem[434] = 10'h1d1;
        mem[435] = 10'h294;
        mem[436] = 10'h179;
        mem[437] = 10'h0ae;
        mem[438] = 10'h057;
        mem[439] = 10'h2f7;
        mem[440] = 10'h38a;
        mem[441] = 10'h0b3;
        mem[442] = 10'h098;
        mem[443] = 10'h31a;
        mem[444] = 10'h2b9;
        mem[445] = 10'h03c;
        mem[446] = 10'h2e2;
        mem[447] = 10'h2ad;
        mem[448] = 10'h170;
        mem[449] = 10'h108;
        mem[450] = 10'h37f;
        mem[451] = 10'h203;
        mem[452] = 10'h129;
        mem[453] = 10'h0a9;
        mem[454] = 10'h3a7;
        mem[455] = 10'h3aa;
        mem[456] = 10'h25e;
        mem[457] = 10'h09f;
        mem[458] = 10'h372;
        mem[459] = 10'h009;
        mem[460] = 10'h24e;
        mem[461] = 10'h1a0;
        mem[462] = 10'h260;
        mem[463] = 10'h0db;
        mem[464] = 10'h024;
        mem[465] = 10'h1a9;
        mem[466] = 10'h110;
        mem[467] = 10'h232;
        mem[468] = 10'h001;
        mem[469] = 10'h3f7;
        mem[470] = 10'h0fa;
        mem[471] = 10'h1cd;
        mem[472] = 10'h22f;
        mem[473] = 10'h0d5;
        mem[474] = 10'h33d;
        mem[475] = 10'h18b;
        mem[476] = 10'h20b;
        mem[477] = 10'h196;
        mem[478] = 10'h0ad;
        mem[479] = 10'h116;
        mem[480] = 10'h2f0;
        mem[481] = 10'h277;
        mem[482] = 10'h2de;
        mem[483] = 10'h04c;
        mem[484] = 10'h17a;
        mem[485] = 10'h2cd;
        mem[486] = 10'h3c4;
        mem[487] = 10'h27d;
        mem[488] = 10'h1d9;
        mem[489] = 10'h02b;
        mem[490] = 10'h3a0;
        mem[491] = 10'h05f;
        mem[492] = 10'h33b;
        mem[493] = 10'h0bb;
        mem[494] = 10'h2db;
        mem[495] = 10'h296;
        mem[496] = 10'h230;
        mem[497] = 10'h3d8;
        mem[498] = 10'h038;
        mem[499] = 10'h12f;
        mem[500] = 10'h295;
        mem[501] = 10'h3a2;
        mem[502] = 10'h151;
        mem[503] = 10'h356;
        mem[504] = 10'h007;
        mem[505] = 10'h267;
        mem[506] = 10'h056;
        mem[507] = 10'h16c;
        mem[508] = 10'h324;
        mem[509] = 10'h0c0;
        mem[510] = 10'h3b0;
        mem[511] = 10'h3c1;
        mem[512] = 10'h3b6;
        mem[513] = 10'h2a7;
        mem[514] = 10'h3b8;
        mem[515] = 10'h09d;
        mem[516] = 10'h0a5;
        mem[517] = 10'h181;
        mem[518] = 10'h3dd;
        mem[519] = 10'h395;
        mem[520] = 10'h1d8;
        mem[521] = 10'h216;
        mem[522] = 10'h191;
        mem[523] = 10'h08e;
        mem[524] = 10'h367;
        mem[525] = 10'h314;
        mem[526] = 10'h313;
        mem[527] = 10'h26b;
        mem[528] = 10'h2c4;
        mem[529] = 10'h1a1;
        mem[530] = 10'h163;
        mem[531] = 10'h23b;
        mem[532] = 10'h289;
        mem[533] = 10'h0a0;
        mem[534] = 10'h025;
        mem[535] = 10'h030;
        mem[536] = 10'h22b;
        mem[537] = 10'h0fe;
        mem[538] = 10'h3b5;
        mem[539] = 10'h3c8;
        mem[540] = 10'h193;
        mem[541] = 10'h301;
        mem[542] = 10'h15e;
        mem[543] = 10'h2ac;
        mem[544] = 10'h0f4;
        mem[545] = 10'h0f9;
        mem[546] = 10'h133;
        mem[547] = 10'h23f;
        mem[548] = 10'h274;
        mem[549] = 10'h37c;
        mem[550] = 10'h3cf;
        mem[551] = 10'h2dd;
        mem[552] = 10'h059;
        mem[553] = 10'h183;
        mem[554] = 10'h097;
        mem[555] = 10'h1cb;
        mem[556] = 10'h1f0;
        mem[557] = 10'h101;
        mem[558] = 10'h206;
        mem[559] = 10'h39d;
        mem[560] = 10'h00c;
        mem[561] = 10'h347;
        mem[562] = 10'h0ec;
        mem[563] = 10'h0ba;
        mem[564] = 10'h080;
        mem[565] = 10'h257;
        mem[566] = 10'h089;
        mem[567] = 10'h17c;
        mem[568] = 10'h2bb;
        mem[569] = 10'h3d6;
        mem[570] = 10'h365;
        mem[571] = 10'h0bd;
        mem[572] = 10'h1e2;
        mem[573] = 10'h1ed;
        mem[574] = 10'h258;
        mem[575] = 10'h280;
        mem[576] = 10'h2d1;
        mem[577] = 10'h1b5;
        mem[578] = 10'h348;
        mem[579] = 10'h161;
        mem[580] = 10'h05a;
        mem[581] = 10'h126;
        mem[582] = 10'h328;
        mem[583] = 10'h392;
        mem[584] = 10'h3ce;
        mem[585] = 10'h3fa;
        mem[586] = 10'h22a;
        mem[587] = 10'h160;
        mem[588] = 10'h0f7;
        mem[589] = 10'h1f3;
        mem[590] = 10'h167;
        mem[591] = 10'h253;
        mem[592] = 10'h369;
        mem[593] = 10'h3a3;
        mem[594] = 10'h1ea;
        mem[595] = 10'h2c0;
        mem[596] = 10'h3ef;
        mem[597] = 10'h111;
        mem[598] = 10'h290;
        mem[599] = 10'h281;
        mem[600] = 10'h1cf;
        mem[601] = 10'h343;
        mem[602] = 10'h00e;
        mem[603] = 10'h1e3;
        mem[604] = 10'h070;
        mem[605] = 10'h0fc;
        mem[606] = 10'h0c7;
        mem[607] = 10'h078;
        mem[608] = 10'h279;
        mem[609] = 10'h32f;
        mem[610] = 10'h10e;
        mem[611] = 10'h376;
        mem[612] = 10'h06d;
        mem[613] = 10'h3bf;
        mem[614] = 10'h2e0;
        mem[615] = 10'h26e;
        mem[616] = 10'h29f;
        mem[617] = 10'h29d;
        mem[618] = 10'h1c3;
        mem[619] = 10'h0af;
        mem[620] = 10'h0b9;
        mem[621] = 10'h14b;
        mem[622] = 10'h11f;
        mem[623] = 10'h020;
        mem[624] = 10'h1e9;
        mem[625] = 10'h164;
        mem[626] = 10'h375;
        mem[627] = 10'h1bd;
        mem[628] = 10'h19c;
        mem[629] = 10'h185;
        mem[630] = 10'h389;
        mem[631] = 10'h2a3;
        mem[632] = 10'h3e1;
        mem[633] = 10'h1f6;
        mem[634] = 10'h1d0;
        mem[635] = 10'h131;
        mem[636] = 10'h12c;
        mem[637] = 10'h022;
        mem[638] = 10'h169;
        mem[639] = 10'h2eb;
        mem[640] = 10'h1c8;
        mem[641] = 10'h2e1;
        mem[642] = 10'h2a5;
        mem[643] = 10'h1ca;
        mem[644] = 10'h0ed;
        mem[645] = 10'h2e6;
        mem[646] = 10'h09a;
        mem[647] = 10'h12a;
        mem[648] = 10'h2ce;
        mem[649] = 10'h27f;
        mem[650] = 10'h318;
        mem[651] = 10'h087;
        mem[652] = 10'h25a;
        mem[653] = 10'h0c5;
        mem[654] = 10'h37b;
        mem[655] = 10'h182;
        mem[656] = 10'h067;
        mem[657] = 10'h040;
        mem[658] = 10'h0f0;
        mem[659] = 10'h379;
        mem[660] = 10'h3ab;
        mem[661] = 10'h0a4;
        mem[662] = 10'h357;
        mem[663] = 10'h1ff;
        mem[664] = 10'h0e8;
        mem[665] = 10'h0d4;
        mem[666] = 10'h008;
        mem[667] = 10'h054;
        mem[668] = 10'h095;
        mem[669] = 10'h340;
        mem[670] = 10'h01f;
        mem[671] = 10'h115;
        mem[672] = 10'h320;
        mem[673] = 10'h1fe;
        mem[674] = 10'h2f5;
        mem[675] = 10'h235;
        mem[676] = 10'h2b4;
        mem[677] = 10'h0a7;
        mem[678] = 10'h159;
        mem[679] = 10'h1a6;
        mem[680] = 10'h0df;
        mem[681] = 10'h157;
        mem[682] = 10'h2e5;
        mem[683] = 10'h252;
        mem[684] = 10'h174;
        mem[685] = 10'h304;
        mem[686] = 10'h11d;
        mem[687] = 10'h000;
        mem[688] = 10'h220;
        mem[689] = 10'h386;
        mem[690] = 10'h30b;
        mem[691] = 10'h2d3;
        mem[692] = 10'h28d;
        mem[693] = 10'h14f;
        mem[694] = 10'h3ed;
        mem[695] = 10'h02c;
        mem[696] = 10'h2ed;
        mem[697] = 10'h130;
        mem[698] = 10'h228;
        mem[699] = 10'h07b;
        mem[700] = 10'h396;
        mem[701] = 10'h0cd;
        mem[702] = 10'h0e2;
        mem[703] = 10'h1ba;
        mem[704] = 10'h394;
        mem[705] = 10'h2b3;
        mem[706] = 10'h1a7;
        mem[707] = 10'h0c8;
        mem[708] = 10'h1a3;
        mem[709] = 10'h16d;
        mem[710] = 10'h2ff;
        mem[711] = 10'h05c;
        mem[712] = 10'h219;
        mem[713] = 10'h3eb;
        mem[714] = 10'h0ab;
        mem[715] = 10'h316;
        mem[716] = 10'h122;
        mem[717] = 10'h0a6;
        mem[718] = 10'h308;
        mem[719] = 10'h109;
        mem[720] = 10'h248;
        mem[721] = 10'h2a6;
        mem[722] = 10'h1b3;
        mem[723] = 10'h205;
        mem[724] = 10'h072;
        mem[725] = 10'h172;
        mem[726] = 10'h005;
        mem[727] = 10'h156;
        mem[728] = 10'h35d;
        mem[729] = 10'h3bc;
        mem[730] = 10'h19d;
        mem[731] = 10'h12e;
        mem[732] = 10'h09c;
        mem[733] = 10'h2ab;
        mem[734] = 10'h346;
        mem[735] = 10'h3e4;
        mem[736] = 10'h0c3;
        mem[737] = 10'h195;
        mem[738] = 10'h01a;
        mem[739] = 10'h238;
        mem[740] = 10'h050;
        mem[741] = 10'h29c;
        mem[742] = 10'h391;
        mem[743] = 10'h031;
        mem[744] = 10'h2a8;
        mem[745] = 10'h01d;
        mem[746] = 10'h2fa;
        mem[747] = 10'h0d9;
        mem[748] = 10'h08d;
        mem[749] = 10'h086;
        mem[750] = 10'h065;
        mem[751] = 10'h075;
        mem[752] = 10'h153;
        mem[753] = 10'h088;
        mem[754] = 10'h021;
        mem[755] = 10'h1a8;
        mem[756] = 10'h377;
        mem[757] = 10'h1fb;
        mem[758] = 10'h3ae;
        mem[759] = 10'h382;
        mem[760] = 10'h13d;
        mem[761] = 10'h11c;
        mem[762] = 10'h158;
        mem[763] = 10'h387;
        mem[764] = 10'h1df;
        mem[765] = 10'h33c;
        mem[766] = 10'h1ac;
        mem[767] = 10'h134;
        mem[768] = 10'h3e9;
        mem[769] = 10'h036;
        mem[770] = 10'h3e2;
        mem[771] = 10'h325;
        mem[772] = 10'h015;
        mem[773] = 10'h1b9;
        mem[774] = 10'h26a;
        mem[775] = 10'h312;
        mem[776] = 10'h0b0;
        mem[777] = 10'h298;
        mem[778] = 10'h0b6;
        mem[779] = 10'h18f;
        mem[780] = 10'h2d2;
        mem[781] = 10'h2e9;
        mem[782] = 10'h35c;
        mem[783] = 10'h284;
        mem[784] = 10'h051;
        mem[785] = 10'h1eb;
        mem[786] = 10'h0b7;
        mem[787] = 10'h28b;
        mem[788] = 10'h210;
        mem[789] = 10'h227;
        mem[790] = 10'h04f;
        mem[791] = 10'h31f;
        mem[792] = 10'h1bf;
        mem[793] = 10'h0eb;
        mem[794] = 10'h326;
        mem[795] = 10'h20c;
        mem[796] = 10'h175;
        mem[797] = 10'h30a;
        mem[798] = 10'h1e7;
        mem[799] = 10'h3df;
        mem[800] = 10'h04a;
        mem[801] = 10'h34b;
        mem[802] = 10'h2f6;
        mem[803] = 10'h241;
        mem[804] = 10'h1a4;
        mem[805] = 10'h202;
        mem[806] = 10'h3a1;
        mem[807] = 10'h1da;
        mem[808] = 10'h19a;
        mem[809] = 10'h06a;
        mem[810] = 10'h35f;
        mem[811] = 10'h32e;
        mem[812] = 10'h068;
        mem[813] = 10'h154;
        mem[814] = 10'h150;
        mem[815] = 10'h01e;
        mem[816] = 10'h184;
        mem[817] = 10'h3bb;
        mem[818] = 10'h1ab;
        mem[819] = 10'h233;
        mem[820] = 10'h0ee;
        mem[821] = 10'h2ba;
        mem[822] = 10'h0b8;
        mem[823] = 10'h079;
        mem[824] = 10'h3cb;
        mem[825] = 10'h18c;
        mem[826] = 10'h1f7;
        mem[827] = 10'h334;
        mem[828] = 10'h00b;
        mem[829] = 10'h1b2;
        mem[830] = 10'h21f;
        mem[831] = 10'h137;
        mem[832] = 10'h187;
        mem[833] = 10'h3e0;
        mem[834] = 10'h276;
        mem[835] = 10'h214;
        mem[836] = 10'h207;
        mem[837] = 10'h2cb;
        mem[838] = 10'h16b;
        mem[839] = 10'h25c;
        mem[840] = 10'h2a4;
        mem[841] = 10'h38e;
        mem[842] = 10'h32a;
        mem[843] = 10'h0c9;
        mem[844] = 10'h123;
        mem[845] = 10'h0b2;
        mem[846] = 10'h128;
        mem[847] = 10'h2bd;
        mem[848] = 10'h29b;
        mem[849] = 10'h125;
        mem[850] = 10'h1c5;
        mem[851] = 10'h3e5;
        mem[852] = 10'h1d2;
        mem[853] = 10'h21d;
        mem[854] = 10'h39e;
        mem[855] = 10'h1b0;
        mem[856] = 10'h3b4;
        mem[857] = 10'h2d7;
        mem[858] = 10'h22e;
        mem[859] = 10'h152;
        mem[860] = 10'h15f;
        mem[861] = 10'h23e;
        mem[862] = 10'h39b;
        mem[863] = 10'h0dc;
        mem[864] = 10'h231;
        mem[865] = 10'h177;
        mem[866] = 10'h085;
        mem[867] = 10'h24a;
        mem[868] = 10'h1f2;
        mem[869] = 10'h026;
        mem[870] = 10'h398;
        mem[871] = 10'h271;
        mem[872] = 10'h2e8;
        mem[873] = 10'h1c2;
        mem[874] = 10'h042;
        mem[875] = 10'h05d;
        mem[876] = 10'h14d;
        mem[877] = 10'h011;
        mem[878] = 10'h2ae;
        mem[879] = 10'h1ef;
        mem[880] = 10'h0cf;
        mem[881] = 10'h2df;
        mem[882] = 10'h30f;
        mem[883] = 10'h1f5;
        mem[884] = 10'h3b9;
        mem[885] = 10'h1c1;
        mem[886] = 10'h12b;
        mem[887] = 10'h1bb;
        mem[888] = 10'h269;
        mem[889] = 10'h186;
        mem[890] = 10'h3a4;
        mem[891] = 10'h22d;
        mem[892] = 10'h14c;
        mem[893] = 10'h3ff;
        mem[894] = 10'h0d0;
        mem[895] = 10'h2c5;
        mem[896] = 10'h2d5;
        mem[897] = 10'h1dd;
        mem[898] = 10'h082;
        mem[899] = 10'h121;
        mem[900] = 10'h1dc;
        mem[901] = 10'h165;
        mem[902] = 10'h3f8;
        mem[903] = 10'h212;
        mem[904] = 10'h18d;
        mem[905] = 10'h192;
        mem[906] = 10'h197;
        mem[907] = 10'h0e3;
        mem[908] = 10'h1e6;
        mem[909] = 10'h1d3;
        mem[910] = 10'h058;
        mem[911] = 10'h166;
        mem[912] = 10'h371;
        mem[913] = 10'h300;
        mem[914] = 10'h24f;
        mem[915] = 10'h2aa;
        mem[916] = 10'h003;
        mem[917] = 10'h3bd;
        mem[918] = 10'h3ad;
        mem[919] = 10'h127;
        mem[920] = 10'h349;
        mem[921] = 10'h10c;
        mem[922] = 10'h149;
        mem[923] = 10'h399;
        mem[924] = 10'h305;
        mem[925] = 10'h26f;
        mem[926] = 10'h1c6;
        mem[927] = 10'h37d;
        mem[928] = 10'h0d1;
        mem[929] = 10'h1ee;
        mem[930] = 10'h39f;
        mem[931] = 10'h0e0;
        mem[932] = 10'h144;
        mem[933] = 10'h3ee;
        mem[934] = 10'h113;
        mem[935] = 10'h381;
        mem[936] = 10'h107;
        mem[937] = 10'h200;
        mem[938] = 10'h0b5;
        mem[939] = 10'h30c;
        mem[940] = 10'h1f4;
        mem[941] = 10'h3ac;
        mem[942] = 10'h0bf;
        mem[943] = 10'h338;
        mem[944] = 10'h3b1;
        mem[945] = 10'h045;
        mem[946] = 10'h08f;
        mem[947] = 10'h3f2;
        mem[948] = 10'h10b;
        mem[949] = 10'h224;
        mem[950] = 10'h32d;
        mem[951] = 10'h1e0;
        mem[952] = 10'h3af;
        mem[953] = 10'h37a;
        mem[954] = 10'h1aa;
        mem[955] = 10'h20d;
        mem[956] = 10'h287;
        mem[957] = 10'h07a;
        mem[958] = 10'h384;
        mem[959] = 10'h331;
        mem[960] = 10'h0cb;
        mem[961] = 10'h2b0;
        mem[962] = 10'h0da;
        mem[963] = 10'h162;
        mem[964] = 10'h1fc;
        mem[965] = 10'h1be;
        mem[966] = 10'h363;
        mem[967] = 10'h012;
        mem[968] = 10'h028;
        mem[969] = 10'h094;
        mem[970] = 10'h292;
        mem[971] = 10'h08a;
        mem[972] = 10'h145;
        mem[973] = 10'h043;
        mem[974] = 10'h29e;
        mem[975] = 10'h02a;
        mem[976] = 10'h0d7;
        mem[977] = 10'h00f;
        mem[978] = 10'h066;
        mem[979] = 10'h17e;
        mem[980] = 10'h118;
        mem[981] = 10'h2fb;
        mem[982] = 10'h0f8;
        mem[983] = 10'h08c;
        mem[984] = 10'h344;
        mem[985] = 10'h3ea;
        mem[986] = 10'h029;
        mem[987] = 10'h1d6;
        mem[988] = 10'h3ec;
        mem[989] = 10'h263;
        mem[990] = 10'h35b;
        mem[991] = 10'h222;
        mem[992] = 10'h1e4;
        mem[993] = 10'h10a;
        mem[994] = 10'h04e;
        mem[995] = 10'h390;
        mem[996] = 10'h317;
        mem[997] = 10'h374;
        mem[998] = 10'h1a5;
        mem[999] = 10'h25b;
        mem[1000] = 10'h302;
        mem[1001] = 10'h360;
        mem[1002] = 10'h132;
        mem[1003] = 10'h2fd;
        mem[1004] = 10'h092;
        mem[1005] = 10'h3c6;
        mem[1006] = 10'h3d9;
        mem[1007] = 10'h3b7;
        mem[1008] = 10'h2ec;
        mem[1009] = 10'h176;
        mem[1010] = 10'h385;
        mem[1011] = 10'h243;
        mem[1012] = 10'h27c;
        mem[1013] = 10'h218;
        mem[1014] = 10'h337;
        mem[1015] = 10'h354;
        mem[1016] = 10'h28f;
        mem[1017] = 10'h3d3;
        mem[1018] = 10'h071;
        mem[1019] = 10'h05b;
        mem[1020] = 10'h189;
        mem[1021] = 10'h247;
        mem[1022] = 10'h0f3;
        mem[1023] = 10'h2af;
    end
endmodule

module odo_sbox_large8(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h37c;
        mem[1] = 10'h3d6;
        mem[2] = 10'h234;
        mem[3] = 10'h166;
        mem[4] = 10'h0bc;
        mem[5] = 10'h0b6;
        mem[6] = 10'h091;
        mem[7] = 10'h2e6;
        mem[8] = 10'h1da;
        mem[9] = 10'h1b8;
        mem[10] = 10'h33f;
        mem[11] = 10'h326;
        mem[12] = 10'h3b0;
        mem[13] = 10'h2a3;
        mem[14] = 10'h3b7;
        mem[15] = 10'h371;
        mem[16] = 10'h17d;
        mem[17] = 10'h31e;
        mem[18] = 10'h301;
        mem[19] = 10'h06b;
        mem[20] = 10'h121;
        mem[21] = 10'h303;
        mem[22] = 10'h0c4;
        mem[23] = 10'h00d;
        mem[24] = 10'h182;
        mem[25] = 10'h253;
        mem[26] = 10'h077;
        mem[27] = 10'h1c0;
        mem[28] = 10'h292;
        mem[29] = 10'h3d2;
        mem[30] = 10'h102;
        mem[31] = 10'h0a3;
        mem[32] = 10'h2d2;
        mem[33] = 10'h30d;
        mem[34] = 10'h0a9;
        mem[35] = 10'h2f4;
        mem[36] = 10'h270;
        mem[37] = 10'h181;
        mem[38] = 10'h1a3;
        mem[39] = 10'h03d;
        mem[40] = 10'h207;
        mem[41] = 10'h2c7;
        mem[42] = 10'h282;
        mem[43] = 10'h164;
        mem[44] = 10'h1c3;
        mem[45] = 10'h088;
        mem[46] = 10'h0db;
        mem[47] = 10'h135;
        mem[48] = 10'h3bc;
        mem[49] = 10'h2b6;
        mem[50] = 10'h08a;
        mem[51] = 10'h3d8;
        mem[52] = 10'h22b;
        mem[53] = 10'h3fd;
        mem[54] = 10'h20c;
        mem[55] = 10'h1b1;
        mem[56] = 10'h1b7;
        mem[57] = 10'h006;
        mem[58] = 10'h1c1;
        mem[59] = 10'h092;
        mem[60] = 10'h134;
        mem[61] = 10'h250;
        mem[62] = 10'h2fd;
        mem[63] = 10'h343;
        mem[64] = 10'h025;
        mem[65] = 10'h260;
        mem[66] = 10'h288;
        mem[67] = 10'h05c;
        mem[68] = 10'h230;
        mem[69] = 10'h03a;
        mem[70] = 10'h206;
        mem[71] = 10'h3b3;
        mem[72] = 10'h007;
        mem[73] = 10'h1fb;
        mem[74] = 10'h149;
        mem[75] = 10'h112;
        mem[76] = 10'h0ee;
        mem[77] = 10'h358;
        mem[78] = 10'h075;
        mem[79] = 10'h322;
        mem[80] = 10'h1ea;
        mem[81] = 10'h3c5;
        mem[82] = 10'h3b4;
        mem[83] = 10'h26c;
        mem[84] = 10'h30e;
        mem[85] = 10'h2f7;
        mem[86] = 10'h208;
        mem[87] = 10'h3bf;
        mem[88] = 10'h157;
        mem[89] = 10'h17c;
        mem[90] = 10'h165;
        mem[91] = 10'h29a;
        mem[92] = 10'h074;
        mem[93] = 10'h2a0;
        mem[94] = 10'h2d0;
        mem[95] = 10'h33a;
        mem[96] = 10'h267;
        mem[97] = 10'h2e5;
        mem[98] = 10'h2ce;
        mem[99] = 10'h251;
        mem[100] = 10'h26a;
        mem[101] = 10'h12d;
        mem[102] = 10'h00e;
        mem[103] = 10'h24f;
        mem[104] = 10'h246;
        mem[105] = 10'h2e4;
        mem[106] = 10'h016;
        mem[107] = 10'h2b2;
        mem[108] = 10'h1be;
        mem[109] = 10'h1eb;
        mem[110] = 10'h190;
        mem[111] = 10'h0e0;
        mem[112] = 10'h078;
        mem[113] = 10'h017;
        mem[114] = 10'h258;
        mem[115] = 10'h1a8;
        mem[116] = 10'h3cb;
        mem[117] = 10'h349;
        mem[118] = 10'h173;
        mem[119] = 10'h0fc;
        mem[120] = 10'h3f2;
        mem[121] = 10'h3df;
        mem[122] = 10'h275;
        mem[123] = 10'h0b7;
        mem[124] = 10'h32e;
        mem[125] = 10'h213;
        mem[126] = 10'h3fe;
        mem[127] = 10'h1ba;
        mem[128] = 10'h045;
        mem[129] = 10'h300;
        mem[130] = 10'h2e9;
        mem[131] = 10'h2f0;
        mem[132] = 10'h191;
        mem[133] = 10'h2dd;
        mem[134] = 10'h07b;
        mem[135] = 10'h1f4;
        mem[136] = 10'h001;
        mem[137] = 10'h3ff;
        mem[138] = 10'h295;
        mem[139] = 10'h080;
        mem[140] = 10'h0ff;
        mem[141] = 10'h348;
        mem[142] = 10'h39c;
        mem[143] = 10'h18c;
        mem[144] = 10'h2a1;
        mem[145] = 10'h02e;
        mem[146] = 10'h353;
        mem[147] = 10'h0ed;
        mem[148] = 10'h27f;
        mem[149] = 10'h2f3;
        mem[150] = 10'h36b;
        mem[151] = 10'h2b7;
        mem[152] = 10'h15e;
        mem[153] = 10'h07f;
        mem[154] = 10'h38d;
        mem[155] = 10'h175;
        mem[156] = 10'h244;
        mem[157] = 10'h3f8;
        mem[158] = 10'h2b9;
        mem[159] = 10'h2c2;
        mem[160] = 10'h18a;
        mem[161] = 10'h2ae;
        mem[162] = 10'h344;
        mem[163] = 10'h08c;
        mem[164] = 10'h08f;
        mem[165] = 10'h2e0;
        mem[166] = 10'h39a;
        mem[167] = 10'h04b;
        mem[168] = 10'h000;
        mem[169] = 10'h043;
        mem[170] = 10'h196;
        mem[171] = 10'h313;
        mem[172] = 10'h105;
        mem[173] = 10'h280;
        mem[174] = 10'h066;
        mem[175] = 10'h171;
        mem[176] = 10'h142;
        mem[177] = 10'h115;
        mem[178] = 10'h312;
        mem[179] = 10'h1f8;
        mem[180] = 10'h1c4;
        mem[181] = 10'h35e;
        mem[182] = 10'h1d2;
        mem[183] = 10'h2d5;
        mem[184] = 10'h29f;
        mem[185] = 10'h0dd;
        mem[186] = 10'h106;
        mem[187] = 10'h194;
        mem[188] = 10'h02c;
        mem[189] = 10'h0a2;
        mem[190] = 10'h068;
        mem[191] = 10'h0da;
        mem[192] = 10'h0bd;
        mem[193] = 10'h221;
        mem[194] = 10'h228;
        mem[195] = 10'h333;
        mem[196] = 10'h396;
        mem[197] = 10'h125;
        mem[198] = 10'h2d9;
        mem[199] = 10'h223;
        mem[200] = 10'h13d;
        mem[201] = 10'h0ab;
        mem[202] = 10'h3de;
        mem[203] = 10'h1e6;
        mem[204] = 10'h202;
        mem[205] = 10'h2bc;
        mem[206] = 10'h394;
        mem[207] = 10'h1ac;
        mem[208] = 10'h08b;
        mem[209] = 10'h19e;
        mem[210] = 10'h1e8;
        mem[211] = 10'h10e;
        mem[212] = 10'h1ae;
        mem[213] = 10'h17a;
        mem[214] = 10'h23f;
        mem[215] = 10'h37f;
        mem[216] = 10'h063;
        mem[217] = 10'h071;
        mem[218] = 10'h318;
        mem[219] = 10'h0cb;
        mem[220] = 10'h369;
        mem[221] = 10'h16f;
        mem[222] = 10'h33b;
        mem[223] = 10'h10d;
        mem[224] = 10'h305;
        mem[225] = 10'h238;
        mem[226] = 10'h252;
        mem[227] = 10'h01a;
        mem[228] = 10'h3ef;
        mem[229] = 10'h12e;
        mem[230] = 10'h17f;
        mem[231] = 10'h19a;
        mem[232] = 10'h1ca;
        mem[233] = 10'h0c3;
        mem[234] = 10'h1d0;
        mem[235] = 10'h031;
        mem[236] = 10'h179;
        mem[237] = 10'h0a5;
        mem[238] = 10'h2c9;
        mem[239] = 10'h33e;
        mem[240] = 10'h29d;
        mem[241] = 10'h085;
        mem[242] = 10'h2cd;
        mem[243] = 10'h1db;
        mem[244] = 10'h220;
        mem[245] = 10'h06e;
        mem[246] = 10'h0f1;
        mem[247] = 10'h23a;
        mem[248] = 10'h3a0;
        mem[249] = 10'h14b;
        mem[250] = 10'h097;
        mem[251] = 10'h231;
        mem[252] = 10'h08e;
        mem[253] = 10'h201;
        mem[254] = 10'h2a5;
        mem[255] = 10'h21f;
        mem[256] = 10'h028;
        mem[257] = 10'h003;
        mem[258] = 10'h1c8;
        mem[259] = 10'h399;
        mem[260] = 10'h024;
        mem[261] = 10'h2ab;
        mem[262] = 10'h3eb;
        mem[263] = 10'h3ae;
        mem[264] = 10'h36f;
        mem[265] = 10'h34b;
        mem[266] = 10'h21c;
        mem[267] = 10'h05f;
        mem[268] = 10'h053;
        mem[269] = 10'h0f9;
        mem[270] = 10'h3bd;
        mem[271] = 10'h082;
        mem[272] = 10'h02d;
        mem[273] = 10'h1a2;
        mem[274] = 10'h224;
        mem[275] = 10'h227;
        mem[276] = 10'h27a;
        mem[277] = 10'h0e7;
        mem[278] = 10'h013;
        mem[279] = 10'h09e;
        mem[280] = 10'h25c;
        mem[281] = 10'h151;
        mem[282] = 10'h055;
        mem[283] = 10'h0e8;
        mem[284] = 10'h347;
        mem[285] = 10'h38a;
        mem[286] = 10'h0c0;
        mem[287] = 10'h20b;
        mem[288] = 10'h393;
        mem[289] = 10'h0e5;
        mem[290] = 10'h033;
        mem[291] = 10'h1e3;
        mem[292] = 10'h07c;
        mem[293] = 10'h242;
        mem[294] = 10'h098;
        mem[295] = 10'h1ee;
        mem[296] = 10'h038;
        mem[297] = 10'h009;
        mem[298] = 10'h375;
        mem[299] = 10'h276;
        mem[300] = 10'h28a;
        mem[301] = 10'h11e;
        mem[302] = 10'h0fe;
        mem[303] = 10'h123;
        mem[304] = 10'h0f0;
        mem[305] = 10'h1aa;
        mem[306] = 10'h10a;
        mem[307] = 10'h189;
        mem[308] = 10'h0ea;
        mem[309] = 10'h39e;
        mem[310] = 10'h047;
        mem[311] = 10'h2a7;
        mem[312] = 10'h19d;
        mem[313] = 10'h31c;
        mem[314] = 10'h3e0;
        mem[315] = 10'h397;
        mem[316] = 10'h114;
        mem[317] = 10'h3ac;
        mem[318] = 10'h0f2;
        mem[319] = 10'h28b;
        mem[320] = 10'h0b2;
        mem[321] = 10'h131;
        mem[322] = 10'h2b1;
        mem[323] = 10'h184;
        mem[324] = 10'h380;
        mem[325] = 10'h1d6;
        mem[326] = 10'h004;
        mem[327] = 10'h0fd;
        mem[328] = 10'h1f2;
        mem[329] = 10'h374;
        mem[330] = 10'h2ac;
        mem[331] = 10'h286;
        mem[332] = 10'h3af;
        mem[333] = 10'h159;
        mem[334] = 10'h0af;
        mem[335] = 10'h081;
        mem[336] = 10'h3c0;
        mem[337] = 10'h15b;
        mem[338] = 10'h1b2;
        mem[339] = 10'h1b6;
        mem[340] = 10'h0de;
        mem[341] = 10'h054;
        mem[342] = 10'h24c;
        mem[343] = 10'h3ea;
        mem[344] = 10'h3ba;
        mem[345] = 10'h1bc;
        mem[346] = 10'h219;
        mem[347] = 10'h0fb;
        mem[348] = 10'h16a;
        mem[349] = 10'h3dc;
        mem[350] = 10'h01d;
        mem[351] = 10'h18e;
        mem[352] = 10'h1af;
        mem[353] = 10'h192;
        mem[354] = 10'h291;
        mem[355] = 10'h23b;
        mem[356] = 10'h29b;
        mem[357] = 10'h143;
        mem[358] = 10'h383;
        mem[359] = 10'h13b;
        mem[360] = 10'h129;
        mem[361] = 10'h060;
        mem[362] = 10'h1e2;
        mem[363] = 10'h345;
        mem[364] = 10'h398;
        mem[365] = 10'h20d;
        mem[366] = 10'h1a5;
        mem[367] = 10'h187;
        mem[368] = 10'h2e3;
        mem[369] = 10'h0a8;
        mem[370] = 10'h32c;
        mem[371] = 10'h372;
        mem[372] = 10'h3da;
        mem[373] = 10'h160;
        mem[374] = 10'h3c1;
        mem[375] = 10'h04a;
        mem[376] = 10'h0ad;
        mem[377] = 10'h2a8;
        mem[378] = 10'h1dd;
        mem[379] = 10'h1f3;
        mem[380] = 10'h1ff;
        mem[381] = 10'h0fa;
        mem[382] = 10'h239;
        mem[383] = 10'h002;
        mem[384] = 10'h3a6;
        mem[385] = 10'h16e;
        mem[386] = 10'h0b1;
        mem[387] = 10'h0c8;
        mem[388] = 10'h156;
        mem[389] = 10'h2ca;
        mem[390] = 10'h340;
        mem[391] = 10'h076;
        mem[392] = 10'h11c;
        mem[393] = 10'h356;
        mem[394] = 10'h2fa;
        mem[395] = 10'h1cc;
        mem[396] = 10'h235;
        mem[397] = 10'h395;
        mem[398] = 10'h36d;
        mem[399] = 10'h061;
        mem[400] = 10'h3d9;
        mem[401] = 10'h1f6;
        mem[402] = 10'h385;
        mem[403] = 10'h1d3;
        mem[404] = 10'h2b8;
        mem[405] = 10'h271;
        mem[406] = 10'h370;
        mem[407] = 10'h34a;
        mem[408] = 10'h1f0;
        mem[409] = 10'h2e8;
        mem[410] = 10'h0bb;
        mem[411] = 10'h128;
        mem[412] = 10'h1e9;
        mem[413] = 10'h176;
        mem[414] = 10'h265;
        mem[415] = 10'h2a6;
        mem[416] = 10'h03f;
        mem[417] = 10'h094;
        mem[418] = 10'h0ce;
        mem[419] = 10'h168;
        mem[420] = 10'h3ad;
        mem[421] = 10'h11f;
        mem[422] = 10'h0d9;
        mem[423] = 10'h109;
        mem[424] = 10'h0e6;
        mem[425] = 10'h0d1;
        mem[426] = 10'h023;
        mem[427] = 10'h214;
        mem[428] = 10'h1a1;
        mem[429] = 10'h20f;
        mem[430] = 10'h243;
        mem[431] = 10'h273;
        mem[432] = 10'h1cb;
        mem[433] = 10'h200;
        mem[434] = 10'h329;
        mem[435] = 10'h2b0;
        mem[436] = 10'h150;
        mem[437] = 10'h3a5;
        mem[438] = 10'h04e;
        mem[439] = 10'h2ee;
        mem[440] = 10'h205;
        mem[441] = 10'h25d;
        mem[442] = 10'h1b0;
        mem[443] = 10'h3f4;
        mem[444] = 10'h26b;
        mem[445] = 10'h14f;
        mem[446] = 10'h2f8;
        mem[447] = 10'h12a;
        mem[448] = 10'h037;
        mem[449] = 10'h064;
        mem[450] = 10'h14a;
        mem[451] = 10'h297;
        mem[452] = 10'h01f;
        mem[453] = 10'h1c9;
        mem[454] = 10'h24e;
        mem[455] = 10'h01e;
        mem[456] = 10'h185;
        mem[457] = 10'h2ba;
        mem[458] = 10'h391;
        mem[459] = 10'h25a;
        mem[460] = 10'h1fa;
        mem[461] = 10'h1d5;
        mem[462] = 10'h14e;
        mem[463] = 10'h320;
        mem[464] = 10'h041;
        mem[465] = 10'h11b;
        mem[466] = 10'h29c;
        mem[467] = 10'h21a;
        mem[468] = 10'h199;
        mem[469] = 10'h2c5;
        mem[470] = 10'h111;
        mem[471] = 10'h018;
        mem[472] = 10'h169;
        mem[473] = 10'h15a;
        mem[474] = 10'h308;
        mem[475] = 10'h3c2;
        mem[476] = 10'h0b5;
        mem[477] = 10'h23c;
        mem[478] = 10'h376;
        mem[479] = 10'h316;
        mem[480] = 10'h13c;
        mem[481] = 10'h28d;
        mem[482] = 10'h00f;
        mem[483] = 10'h384;
        mem[484] = 10'h09b;
        mem[485] = 10'h090;
        mem[486] = 10'h1ec;
        mem[487] = 10'h3b8;
        mem[488] = 10'h22e;
        mem[489] = 10'h390;
        mem[490] = 10'h03e;
        mem[491] = 10'h153;
        mem[492] = 10'h177;
        mem[493] = 10'h257;
        mem[494] = 10'h05a;
        mem[495] = 10'h048;
        mem[496] = 10'h130;
        mem[497] = 10'h0be;
        mem[498] = 10'h1e4;
        mem[499] = 10'h13f;
        mem[500] = 10'h16c;
        mem[501] = 10'h330;
        mem[502] = 10'h17e;
        mem[503] = 10'h3cf;
        mem[504] = 10'h3f5;
        mem[505] = 10'h39f;
        mem[506] = 10'h22c;
        mem[507] = 10'h284;
        mem[508] = 10'h093;
        mem[509] = 10'h212;
        mem[510] = 10'h266;
        mem[511] = 10'h3a7;
        mem[512] = 10'h127;
        mem[513] = 10'h29e;
        mem[514] = 10'h366;
        mem[515] = 10'h331;
        mem[516] = 10'h259;
        mem[517] = 10'h210;
        mem[518] = 10'h27e;
        mem[519] = 10'h116;
        mem[520] = 10'h1a7;
        mem[521] = 10'h324;
        mem[522] = 10'h1de;
        mem[523] = 10'h306;
        mem[524] = 10'h0f8;
        mem[525] = 10'h28c;
        mem[526] = 10'h1b9;
        mem[527] = 10'h139;
        mem[528] = 10'h25f;
        mem[529] = 10'h10c;
        mem[530] = 10'h022;
        mem[531] = 10'h2cc;
        mem[532] = 10'h170;
        mem[533] = 10'h14c;
        mem[534] = 10'h3fc;
        mem[535] = 10'h058;
        mem[536] = 10'h325;
        mem[537] = 10'h3d0;
        mem[538] = 10'h161;
        mem[539] = 10'h0b8;
        mem[540] = 10'h1c5;
        mem[541] = 10'h0df;
        mem[542] = 10'h38c;
        mem[543] = 10'h30f;
        mem[544] = 10'h0cc;
        mem[545] = 10'h3f0;
        mem[546] = 10'h31a;
        mem[547] = 10'h3db;
        mem[548] = 10'h1cf;
        mem[549] = 10'h3c7;
        mem[550] = 10'h0cd;
        mem[551] = 10'h036;
        mem[552] = 10'h3aa;
        mem[553] = 10'h039;
        mem[554] = 10'h141;
        mem[555] = 10'h0d8;
        mem[556] = 10'h334;
        mem[557] = 10'h31b;
        mem[558] = 10'h005;
        mem[559] = 10'h28e;
        mem[560] = 10'h25e;
        mem[561] = 10'h373;
        mem[562] = 10'h070;
        mem[563] = 10'h15c;
        mem[564] = 10'h174;
        mem[565] = 10'h2db;
        mem[566] = 10'h12c;
        mem[567] = 10'h290;
        mem[568] = 10'h26d;
        mem[569] = 10'h140;
        mem[570] = 10'h1d1;
        mem[571] = 10'h215;
        mem[572] = 10'h193;
        mem[573] = 10'h35d;
        mem[574] = 10'h152;
        mem[575] = 10'h22f;
        mem[576] = 10'h087;
        mem[577] = 10'h30a;
        mem[578] = 10'h350;
        mem[579] = 10'h124;
        mem[580] = 10'h3e8;
        mem[581] = 10'h32a;
        mem[582] = 10'h294;
        mem[583] = 10'h0e3;
        mem[584] = 10'h363;
        mem[585] = 10'h3f1;
        mem[586] = 10'h0a0;
        mem[587] = 10'h1f1;
        mem[588] = 10'h1dc;
        mem[589] = 10'h3ec;
        mem[590] = 10'h354;
        mem[591] = 10'h351;
        mem[592] = 10'h132;
        mem[593] = 10'h274;
        mem[594] = 10'h059;
        mem[595] = 10'h0ef;
        mem[596] = 10'h137;
        mem[597] = 10'h3f3;
        mem[598] = 10'h23d;
        mem[599] = 10'h034;
        mem[600] = 10'h03c;
        mem[601] = 10'h15f;
        mem[602] = 10'h079;
        mem[603] = 10'h37e;
        mem[604] = 10'h0cf;
        mem[605] = 10'h30c;
        mem[606] = 10'h015;
        mem[607] = 10'h247;
        mem[608] = 10'h0ae;
        mem[609] = 10'h07e;
        mem[610] = 10'h3e6;
        mem[611] = 10'h2d4;
        mem[612] = 10'h16d;
        mem[613] = 10'h1d4;
        mem[614] = 10'h2ea;
        mem[615] = 10'h3a8;
        mem[616] = 10'h277;
        mem[617] = 10'h1f9;
        mem[618] = 10'h18d;
        mem[619] = 10'h381;
        mem[620] = 10'h183;
        mem[621] = 10'h052;
        mem[622] = 10'h04f;
        mem[623] = 10'h3c8;
        mem[624] = 10'h19f;
        mem[625] = 10'h3c4;
        mem[626] = 10'h0a6;
        mem[627] = 10'h226;
        mem[628] = 10'h0c7;
        mem[629] = 10'h117;
        mem[630] = 10'h3c3;
        mem[631] = 10'h138;
        mem[632] = 10'h0f3;
        mem[633] = 10'h1b5;
        mem[634] = 10'h133;
        mem[635] = 10'h263;
        mem[636] = 10'h245;
        mem[637] = 10'h3a4;
        mem[638] = 10'h248;
        mem[639] = 10'h197;
        mem[640] = 10'h1fc;
        mem[641] = 10'h1fe;
        mem[642] = 10'h0c2;
        mem[643] = 10'h08d;
        mem[644] = 10'h262;
        mem[645] = 10'h09a;
        mem[646] = 10'h104;
        mem[647] = 10'h278;
        mem[648] = 10'h0d3;
        mem[649] = 10'h323;
        mem[650] = 10'h1b4;
        mem[651] = 10'h33c;
        mem[652] = 10'h2de;
        mem[653] = 10'h27c;
        mem[654] = 10'h01b;
        mem[655] = 10'h3ce;
        mem[656] = 10'h040;
        mem[657] = 10'h309;
        mem[658] = 10'h148;
        mem[659] = 10'h20e;
        mem[660] = 10'h3a9;
        mem[661] = 10'h012;
        mem[662] = 10'h35b;
        mem[663] = 10'h3e4;
        mem[664] = 10'h0bf;
        mem[665] = 10'h0e2;
        mem[666] = 10'h34e;
        mem[667] = 10'h3b5;
        mem[668] = 10'h11a;
        mem[669] = 10'h2ff;
        mem[670] = 10'h108;
        mem[671] = 10'h00b;
        mem[672] = 10'h158;
        mem[673] = 10'h178;
        mem[674] = 10'h268;
        mem[675] = 10'h1e7;
        mem[676] = 10'h386;
        mem[677] = 10'h279;
        mem[678] = 10'h307;
        mem[679] = 10'h2d3;
        mem[680] = 10'h362;
        mem[681] = 10'h155;
        mem[682] = 10'h328;
        mem[683] = 10'h232;
        mem[684] = 10'h095;
        mem[685] = 10'h0d7;
        mem[686] = 10'h084;
        mem[687] = 10'h126;
        mem[688] = 10'h21d;
        mem[689] = 10'h3f9;
        mem[690] = 10'h162;
        mem[691] = 10'h056;
        mem[692] = 10'h2f1;
        mem[693] = 10'h365;
        mem[694] = 10'h2e7;
        mem[695] = 10'h1ef;
        mem[696] = 10'h00a;
        mem[697] = 10'h019;
        mem[698] = 10'h073;
        mem[699] = 10'h3b2;
        mem[700] = 10'h086;
        mem[701] = 10'h2dc;
        mem[702] = 10'h0ca;
        mem[703] = 10'h233;
        mem[704] = 10'h269;
        mem[705] = 10'h0b4;
        mem[706] = 10'h3cc;
        mem[707] = 10'h1c6;
        mem[708] = 10'h049;
        mem[709] = 10'h2f6;
        mem[710] = 10'h2df;
        mem[711] = 10'h0f4;
        mem[712] = 10'h057;
        mem[713] = 10'h0d0;
        mem[714] = 10'h1f7;
        mem[715] = 10'h01c;
        mem[716] = 10'h1cd;
        mem[717] = 10'h1c2;
        mem[718] = 10'h3e3;
        mem[719] = 10'h37b;
        mem[720] = 10'h203;
        mem[721] = 10'h180;
        mem[722] = 10'h0c1;
        mem[723] = 10'h1c7;
        mem[724] = 10'h026;
        mem[725] = 10'h332;
        mem[726] = 10'h035;
        mem[727] = 10'h17b;
        mem[728] = 10'h341;
        mem[729] = 10'h07a;
        mem[730] = 10'h209;
        mem[731] = 10'h103;
        mem[732] = 10'h3fa;
        mem[733] = 10'h0eb;
        mem[734] = 10'h37d;
        mem[735] = 10'h0c6;
        mem[736] = 10'h0b0;
        mem[737] = 10'h0f5;
        mem[738] = 10'h032;
        mem[739] = 10'h38e;
        mem[740] = 10'h36a;
        mem[741] = 10'h38f;
        mem[742] = 10'h218;
        mem[743] = 10'h06f;
        mem[744] = 10'h0a4;
        mem[745] = 10'h3b9;
        mem[746] = 10'h147;
        mem[747] = 10'h0d5;
        mem[748] = 10'h337;
        mem[749] = 10'h1e0;
        mem[750] = 10'h367;
        mem[751] = 10'h302;
        mem[752] = 10'h2eb;
        mem[753] = 10'h198;
        mem[754] = 10'h39b;
        mem[755] = 10'h1ab;
        mem[756] = 10'h2cf;
        mem[757] = 10'h225;
        mem[758] = 10'h3fb;
        mem[759] = 10'h3f7;
        mem[760] = 10'h39d;
        mem[761] = 10'h3bb;
        mem[762] = 10'h35f;
        mem[763] = 10'h22d;
        mem[764] = 10'h11d;
        mem[765] = 10'h008;
        mem[766] = 10'h2b4;
        mem[767] = 10'h1b3;
        mem[768] = 10'h067;
        mem[769] = 10'h2f2;
        mem[770] = 10'h0e9;
        mem[771] = 10'h163;
        mem[772] = 10'h14d;
        mem[773] = 10'h2ed;
        mem[774] = 10'h12f;
        mem[775] = 10'h254;
        mem[776] = 10'h2f9;
        mem[777] = 10'h04d;
        mem[778] = 10'h26e;
        mem[779] = 10'h0ec;
        mem[780] = 10'h021;
        mem[781] = 10'h13a;
        mem[782] = 10'h2bf;
        mem[783] = 10'h364;
        mem[784] = 10'h379;
        mem[785] = 10'h027;
        mem[786] = 10'h304;
        mem[787] = 10'h317;
        mem[788] = 10'h2c3;
        mem[789] = 10'h3e1;
        mem[790] = 10'h09f;
        mem[791] = 10'h089;
        mem[792] = 10'h1ad;
        mem[793] = 10'h24d;
        mem[794] = 10'h35a;
        mem[795] = 10'h382;
        mem[796] = 10'h083;
        mem[797] = 10'h2a9;
        mem[798] = 10'h315;
        mem[799] = 10'h2f5;
        mem[800] = 10'h37a;
        mem[801] = 10'h2be;
        mem[802] = 10'h368;
        mem[803] = 10'h186;
        mem[804] = 10'h3ed;
        mem[805] = 10'h222;
        mem[806] = 10'h3d4;
        mem[807] = 10'h34f;
        mem[808] = 10'h0a7;
        mem[809] = 10'h12b;
        mem[810] = 10'h03b;
        mem[811] = 10'h2c0;
        mem[812] = 10'h388;
        mem[813] = 10'h118;
        mem[814] = 10'h261;
        mem[815] = 10'h2ad;
        mem[816] = 10'h030;
        mem[817] = 10'h3cd;
        mem[818] = 10'h119;
        mem[819] = 10'h1fd;
        mem[820] = 10'h00c;
        mem[821] = 10'h359;
        mem[822] = 10'h361;
        mem[823] = 10'h3e5;
        mem[824] = 10'h020;
        mem[825] = 10'h1ce;
        mem[826] = 10'h36c;
        mem[827] = 10'h3a2;
        mem[828] = 10'h249;
        mem[829] = 10'h1e1;
        mem[830] = 10'h1bd;
        mem[831] = 10'h2c6;
        mem[832] = 10'h26f;
        mem[833] = 10'h293;
        mem[834] = 10'h2fc;
        mem[835] = 10'h011;
        mem[836] = 10'h3ca;
        mem[837] = 10'h30b;
        mem[838] = 10'h19b;
        mem[839] = 10'h051;
        mem[840] = 10'h285;
        mem[841] = 10'h0d4;
        mem[842] = 10'h3a1;
        mem[843] = 10'h195;
        mem[844] = 10'h2c8;
        mem[845] = 10'h360;
        mem[846] = 10'h02f;
        mem[847] = 10'h2b5;
        mem[848] = 10'h3c6;
        mem[849] = 10'h0e4;
        mem[850] = 10'h314;
        mem[851] = 10'h069;
        mem[852] = 10'h0e1;
        mem[853] = 10'h3e2;
        mem[854] = 10'h09c;
        mem[855] = 10'h32b;
        mem[856] = 10'h144;
        mem[857] = 10'h3ab;
        mem[858] = 10'h357;
        mem[859] = 10'h029;
        mem[860] = 10'h32d;
        mem[861] = 10'h0aa;
        mem[862] = 10'h0ac;
        mem[863] = 10'h2da;
        mem[864] = 10'h25b;
        mem[865] = 10'h241;
        mem[866] = 10'h28f;
        mem[867] = 10'h18f;
        mem[868] = 10'h2e1;
        mem[869] = 10'h298;
        mem[870] = 10'h0a1;
        mem[871] = 10'h065;
        mem[872] = 10'h1a9;
        mem[873] = 10'h09d;
        mem[874] = 10'h2c1;
        mem[875] = 10'h154;
        mem[876] = 10'h3be;
        mem[877] = 10'h2d1;
        mem[878] = 10'h172;
        mem[879] = 10'h05e;
        mem[880] = 10'h072;
        mem[881] = 10'h311;
        mem[882] = 10'h38b;
        mem[883] = 10'h042;
        mem[884] = 10'h0d2;
        mem[885] = 10'h0f6;
        mem[886] = 10'h3c9;
        mem[887] = 10'h0c9;
        mem[888] = 10'h06c;
        mem[889] = 10'h346;
        mem[890] = 10'h2ef;
        mem[891] = 10'h3d5;
        mem[892] = 10'h3ee;
        mem[893] = 10'h31d;
        mem[894] = 10'h0ba;
        mem[895] = 10'h281;
        mem[896] = 10'h1d8;
        mem[897] = 10'h287;
        mem[898] = 10'h338;
        mem[899] = 10'h1a0;
        mem[900] = 10'h237;
        mem[901] = 10'h04c;
        mem[902] = 10'h335;
        mem[903] = 10'h1bb;
        mem[904] = 10'h283;
        mem[905] = 10'h10b;
        mem[906] = 10'h204;
        mem[907] = 10'h355;
        mem[908] = 10'h336;
        mem[909] = 10'h3b6;
        mem[910] = 10'h2a2;
        mem[911] = 10'h05b;
        mem[912] = 10'h236;
        mem[913] = 10'h06d;
        mem[914] = 10'h34c;
        mem[915] = 10'h3e9;
        mem[916] = 10'h36e;
        mem[917] = 10'h1a6;
        mem[918] = 10'h145;
        mem[919] = 10'h389;
        mem[920] = 10'h2c4;
        mem[921] = 10'h352;
        mem[922] = 10'h02a;
        mem[923] = 10'h229;
        mem[924] = 10'h2fb;
        mem[925] = 10'h310;
        mem[926] = 10'h3a3;
        mem[927] = 10'h21e;
        mem[928] = 10'h378;
        mem[929] = 10'h20a;
        mem[930] = 10'h387;
        mem[931] = 10'h101;
        mem[932] = 10'h31f;
        mem[933] = 10'h010;
        mem[934] = 10'h255;
        mem[935] = 10'h113;
        mem[936] = 10'h2e2;
        mem[937] = 10'h0f7;
        mem[938] = 10'h296;
        mem[939] = 10'h27d;
        mem[940] = 10'h2aa;
        mem[941] = 10'h216;
        mem[942] = 10'h05d;
        mem[943] = 10'h18b;
        mem[944] = 10'h2d8;
        mem[945] = 10'h107;
        mem[946] = 10'h33d;
        mem[947] = 10'h0c5;
        mem[948] = 10'h342;
        mem[949] = 10'h22a;
        mem[950] = 10'h377;
        mem[951] = 10'h3e7;
        mem[952] = 10'h2a4;
        mem[953] = 10'h014;
        mem[954] = 10'h100;
        mem[955] = 10'h2d7;
        mem[956] = 10'h2ec;
        mem[957] = 10'h1e5;
        mem[958] = 10'h06a;
        mem[959] = 10'h044;
        mem[960] = 10'h24b;
        mem[961] = 10'h1bf;
        mem[962] = 10'h10f;
        mem[963] = 10'h2bb;
        mem[964] = 10'h1ed;
        mem[965] = 10'h16b;
        mem[966] = 10'h299;
        mem[967] = 10'h13e;
        mem[968] = 10'h2cb;
        mem[969] = 10'h188;
        mem[970] = 10'h07d;
        mem[971] = 10'h15d;
        mem[972] = 10'h3b1;
        mem[973] = 10'h24a;
        mem[974] = 10'h02b;
        mem[975] = 10'h122;
        mem[976] = 10'h0d6;
        mem[977] = 10'h046;
        mem[978] = 10'h27b;
        mem[979] = 10'h21b;
        mem[980] = 10'h096;
        mem[981] = 10'h2af;
        mem[982] = 10'h0b3;
        mem[983] = 10'h32f;
        mem[984] = 10'h1d9;
        mem[985] = 10'h3d1;
        mem[986] = 10'h392;
        mem[987] = 10'h3d7;
        mem[988] = 10'h19c;
        mem[989] = 10'h110;
        mem[990] = 10'h23e;
        mem[991] = 10'h264;
        mem[992] = 10'h167;
        mem[993] = 10'h1a4;
        mem[994] = 10'h34d;
        mem[995] = 10'h319;
        mem[996] = 10'h0b9;
        mem[997] = 10'h272;
        mem[998] = 10'h062;
        mem[999] = 10'h339;
        mem[1000] = 10'h240;
        mem[1001] = 10'h0dc;
        mem[1002] = 10'h1d7;
        mem[1003] = 10'h35c;
        mem[1004] = 10'h256;
        mem[1005] = 10'h050;
        mem[1006] = 10'h3dd;
        mem[1007] = 10'h2d6;
        mem[1008] = 10'h327;
        mem[1009] = 10'h2bd;
        mem[1010] = 10'h289;
        mem[1011] = 10'h2b3;
        mem[1012] = 10'h211;
        mem[1013] = 10'h3d3;
        mem[1014] = 10'h1f5;
        mem[1015] = 10'h1df;
        mem[1016] = 10'h3f6;
        mem[1017] = 10'h2fe;
        mem[1018] = 10'h099;
        mem[1019] = 10'h217;
        mem[1020] = 10'h120;
        mem[1021] = 10'h321;
        mem[1022] = 10'h146;
        mem[1023] = 10'h136;
    end
endmodule

module odo_sbox_large9(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h2f6;
        mem[1] = 10'h36c;
        mem[2] = 10'h167;
        mem[3] = 10'h226;
        mem[4] = 10'h2c2;
        mem[5] = 10'h22e;
        mem[6] = 10'h03a;
        mem[7] = 10'h308;
        mem[8] = 10'h10a;
        mem[9] = 10'h231;
        mem[10] = 10'h171;
        mem[11] = 10'h3fa;
        mem[12] = 10'h2fd;
        mem[13] = 10'h389;
        mem[14] = 10'h0a0;
        mem[15] = 10'h1e9;
        mem[16] = 10'h2b7;
        mem[17] = 10'h17c;
        mem[18] = 10'h3a9;
        mem[19] = 10'h23b;
        mem[20] = 10'h172;
        mem[21] = 10'h22c;
        mem[22] = 10'h1ca;
        mem[23] = 10'h342;
        mem[24] = 10'h1c3;
        mem[25] = 10'h173;
        mem[26] = 10'h0a5;
        mem[27] = 10'h1bd;
        mem[28] = 10'h0cc;
        mem[29] = 10'h0b6;
        mem[30] = 10'h322;
        mem[31] = 10'h336;
        mem[32] = 10'h209;
        mem[33] = 10'h38f;
        mem[34] = 10'h2c4;
        mem[35] = 10'h0de;
        mem[36] = 10'h32f;
        mem[37] = 10'h208;
        mem[38] = 10'h0f6;
        mem[39] = 10'h1a9;
        mem[40] = 10'h3fc;
        mem[41] = 10'h3d7;
        mem[42] = 10'h1fa;
        mem[43] = 10'h22a;
        mem[44] = 10'h220;
        mem[45] = 10'h2a7;
        mem[46] = 10'h377;
        mem[47] = 10'h17f;
        mem[48] = 10'h29a;
        mem[49] = 10'h3b7;
        mem[50] = 10'h3a1;
        mem[51] = 10'h083;
        mem[52] = 10'h3e5;
        mem[53] = 10'h26b;
        mem[54] = 10'h349;
        mem[55] = 10'h162;
        mem[56] = 10'h3d5;
        mem[57] = 10'h2e7;
        mem[58] = 10'h1a8;
        mem[59] = 10'h16d;
        mem[60] = 10'h163;
        mem[61] = 10'h044;
        mem[62] = 10'h081;
        mem[63] = 10'h0b5;
        mem[64] = 10'h3b0;
        mem[65] = 10'h243;
        mem[66] = 10'h225;
        mem[67] = 10'h2aa;
        mem[68] = 10'h065;
        mem[69] = 10'h3f4;
        mem[70] = 10'h217;
        mem[71] = 10'h066;
        mem[72] = 10'h26a;
        mem[73] = 10'h00b;
        mem[74] = 10'h3f1;
        mem[75] = 10'h01f;
        mem[76] = 10'h004;
        mem[77] = 10'h283;
        mem[78] = 10'h3a7;
        mem[79] = 10'h3e8;
        mem[80] = 10'h15a;
        mem[81] = 10'h024;
        mem[82] = 10'h256;
        mem[83] = 10'h2da;
        mem[84] = 10'h091;
        mem[85] = 10'h1d2;
        mem[86] = 10'h10d;
        mem[87] = 10'h1a6;
        mem[88] = 10'h188;
        mem[89] = 10'h3bf;
        mem[90] = 10'h0a8;
        mem[91] = 10'h268;
        mem[92] = 10'h19d;
        mem[93] = 10'h28a;
        mem[94] = 10'h17a;
        mem[95] = 10'h1ea;
        mem[96] = 10'h2ba;
        mem[97] = 10'h221;
        mem[98] = 10'h1f1;
        mem[99] = 10'h222;
        mem[100] = 10'h272;
        mem[101] = 10'h2a1;
        mem[102] = 10'h045;
        mem[103] = 10'h18c;
        mem[104] = 10'h38c;
        mem[105] = 10'h1df;
        mem[106] = 10'h1cd;
        mem[107] = 10'h183;
        mem[108] = 10'h05c;
        mem[109] = 10'h3f2;
        mem[110] = 10'h12f;
        mem[111] = 10'h3f5;
        mem[112] = 10'h0c7;
        mem[113] = 10'h12a;
        mem[114] = 10'h1b5;
        mem[115] = 10'h3b9;
        mem[116] = 10'h052;
        mem[117] = 10'h2e0;
        mem[118] = 10'h305;
        mem[119] = 10'h064;
        mem[120] = 10'h2dd;
        mem[121] = 10'h2dc;
        mem[122] = 10'h24c;
        mem[123] = 10'h1fe;
        mem[124] = 10'h2ab;
        mem[125] = 10'h20a;
        mem[126] = 10'h242;
        mem[127] = 10'h27a;
        mem[128] = 10'h013;
        mem[129] = 10'h2ff;
        mem[130] = 10'h291;
        mem[131] = 10'h396;
        mem[132] = 10'h310;
        mem[133] = 10'h1e5;
        mem[134] = 10'h355;
        mem[135] = 10'h2c0;
        mem[136] = 10'h195;
        mem[137] = 10'h2ea;
        mem[138] = 10'h1b4;
        mem[139] = 10'h0f2;
        mem[140] = 10'h3ec;
        mem[141] = 10'h043;
        mem[142] = 10'h061;
        mem[143] = 10'h33a;
        mem[144] = 10'h3d9;
        mem[145] = 10'h0c1;
        mem[146] = 10'h3bb;
        mem[147] = 10'h1d9;
        mem[148] = 10'h1e2;
        mem[149] = 10'h2c9;
        mem[150] = 10'h154;
        mem[151] = 10'h14f;
        mem[152] = 10'h384;
        mem[153] = 10'h08d;
        mem[154] = 10'h0eb;
        mem[155] = 10'h0c0;
        mem[156] = 10'h146;
        mem[157] = 10'h1f4;
        mem[158] = 10'h1d1;
        mem[159] = 10'h1ff;
        mem[160] = 10'h143;
        mem[161] = 10'h223;
        mem[162] = 10'h319;
        mem[163] = 10'h3fd;
        mem[164] = 10'h1c8;
        mem[165] = 10'h05f;
        mem[166] = 10'h239;
        mem[167] = 10'h3cc;
        mem[168] = 10'h210;
        mem[169] = 10'h187;
        mem[170] = 10'h01e;
        mem[171] = 10'h2c3;
        mem[172] = 10'h34e;
        mem[173] = 10'h2c5;
        mem[174] = 10'h3a6;
        mem[175] = 10'h3b4;
        mem[176] = 10'h2be;
        mem[177] = 10'h206;
        mem[178] = 10'h1de;
        mem[179] = 10'h1a0;
        mem[180] = 10'h2a9;
        mem[181] = 10'h03e;
        mem[182] = 10'h288;
        mem[183] = 10'h0ec;
        mem[184] = 10'h21a;
        mem[185] = 10'h014;
        mem[186] = 10'h0e9;
        mem[187] = 10'h2ef;
        mem[188] = 10'h3ee;
        mem[189] = 10'h0db;
        mem[190] = 10'h121;
        mem[191] = 10'h278;
        mem[192] = 10'h30c;
        mem[193] = 10'h07c;
        mem[194] = 10'h385;
        mem[195] = 10'h266;
        mem[196] = 10'h304;
        mem[197] = 10'h082;
        mem[198] = 10'h0a7;
        mem[199] = 10'h0d5;
        mem[200] = 10'h0d0;
        mem[201] = 10'h1db;
        mem[202] = 10'h271;
        mem[203] = 10'h330;
        mem[204] = 10'h229;
        mem[205] = 10'h382;
        mem[206] = 10'h1a7;
        mem[207] = 10'h0e3;
        mem[208] = 10'h3cb;
        mem[209] = 10'h11f;
        mem[210] = 10'h113;
        mem[211] = 10'h27f;
        mem[212] = 10'h388;
        mem[213] = 10'h35d;
        mem[214] = 10'h1d6;
        mem[215] = 10'h2d3;
        mem[216] = 10'h0e2;
        mem[217] = 10'h14e;
        mem[218] = 10'h257;
        mem[219] = 10'h3dd;
        mem[220] = 10'h192;
        mem[221] = 10'h366;
        mem[222] = 10'h286;
        mem[223] = 10'h359;
        mem[224] = 10'h2d9;
        mem[225] = 10'h23c;
        mem[226] = 10'h372;
        mem[227] = 10'h32c;
        mem[228] = 10'h3ed;
        mem[229] = 10'h249;
        mem[230] = 10'h380;
        mem[231] = 10'h2b3;
        mem[232] = 10'h18b;
        mem[233] = 10'h29d;
        mem[234] = 10'h392;
        mem[235] = 10'h259;
        mem[236] = 10'h253;
        mem[237] = 10'h3ae;
        mem[238] = 10'h184;
        mem[239] = 10'h275;
        mem[240] = 10'h320;
        mem[241] = 10'h204;
        mem[242] = 10'h152;
        mem[243] = 10'h2eb;
        mem[244] = 10'h092;
        mem[245] = 10'h21e;
        mem[246] = 10'h0ad;
        mem[247] = 10'h3b1;
        mem[248] = 10'h03b;
        mem[249] = 10'h158;
        mem[250] = 10'h3eb;
        mem[251] = 10'h376;
        mem[252] = 10'h258;
        mem[253] = 10'h3de;
        mem[254] = 10'h36a;
        mem[255] = 10'h094;
        mem[256] = 10'h33f;
        mem[257] = 10'h1cc;
        mem[258] = 10'h3cd;
        mem[259] = 10'h27e;
        mem[260] = 10'h247;
        mem[261] = 10'h23d;
        mem[262] = 10'h25d;
        mem[263] = 10'h34b;
        mem[264] = 10'h027;
        mem[265] = 10'h2fb;
        mem[266] = 10'h112;
        mem[267] = 10'h0b4;
        mem[268] = 10'h325;
        mem[269] = 10'h134;
        mem[270] = 10'h35e;
        mem[271] = 10'h1f2;
        mem[272] = 10'h362;
        mem[273] = 10'h090;
        mem[274] = 10'h2e8;
        mem[275] = 10'h02a;
        mem[276] = 10'h07d;
        mem[277] = 10'h26d;
        mem[278] = 10'h150;
        mem[279] = 10'h2a4;
        mem[280] = 10'h387;
        mem[281] = 10'h16b;
        mem[282] = 10'h2d6;
        mem[283] = 10'h022;
        mem[284] = 10'h28f;
        mem[285] = 10'h15c;
        mem[286] = 10'h35f;
        mem[287] = 10'h269;
        mem[288] = 10'h177;
        mem[289] = 10'h14a;
        mem[290] = 10'h0ba;
        mem[291] = 10'h267;
        mem[292] = 10'h057;
        mem[293] = 10'h340;
        mem[294] = 10'h11e;
        mem[295] = 10'h030;
        mem[296] = 10'h30a;
        mem[297] = 10'h1b8;
        mem[298] = 10'h18a;
        mem[299] = 10'h20e;
        mem[300] = 10'h2bf;
        mem[301] = 10'h0a4;
        mem[302] = 10'h373;
        mem[303] = 10'h3c2;
        mem[304] = 10'h13f;
        mem[305] = 10'h1f5;
        mem[306] = 10'h00c;
        mem[307] = 10'h1ee;
        mem[308] = 10'h12e;
        mem[309] = 10'h07a;
        mem[310] = 10'h1f0;
        mem[311] = 10'h292;
        mem[312] = 10'h28b;
        mem[313] = 10'h334;
        mem[314] = 10'h37c;
        mem[315] = 10'h020;
        mem[316] = 10'h120;
        mem[317] = 10'h3e9;
        mem[318] = 10'h10c;
        mem[319] = 10'h3ce;
        mem[320] = 10'h1e1;
        mem[321] = 10'h1f6;
        mem[322] = 10'h0e8;
        mem[323] = 10'h137;
        mem[324] = 10'h393;
        mem[325] = 10'h3ff;
        mem[326] = 10'h0af;
        mem[327] = 10'h2ad;
        mem[328] = 10'h3cf;
        mem[329] = 10'h279;
        mem[330] = 10'h205;
        mem[331] = 10'h034;
        mem[332] = 10'h0ee;
        mem[333] = 10'h26c;
        mem[334] = 10'h0fb;
        mem[335] = 10'h2e4;
        mem[336] = 10'h05b;
        mem[337] = 10'h144;
        mem[338] = 10'h005;
        mem[339] = 10'h105;
        mem[340] = 10'h21b;
        mem[341] = 10'h186;
        mem[342] = 10'h27c;
        mem[343] = 10'h24e;
        mem[344] = 10'h099;
        mem[345] = 10'h04d;
        mem[346] = 10'h0a6;
        mem[347] = 10'h236;
        mem[348] = 10'h3e3;
        mem[349] = 10'h0e6;
        mem[350] = 10'h33d;
        mem[351] = 10'h036;
        mem[352] = 10'h0d7;
        mem[353] = 10'h213;
        mem[354] = 10'h341;
        mem[355] = 10'h159;
        mem[356] = 10'h0be;
        mem[357] = 10'h15f;
        mem[358] = 10'h32b;
        mem[359] = 10'h124;
        mem[360] = 10'h285;
        mem[361] = 10'h2d8;
        mem[362] = 10'h297;
        mem[363] = 10'h273;
        mem[364] = 10'h3d4;
        mem[365] = 10'h0ae;
        mem[366] = 10'h3f3;
        mem[367] = 10'h26f;
        mem[368] = 10'h2f8;
        mem[369] = 10'h346;
        mem[370] = 10'h106;
        mem[371] = 10'h300;
        mem[372] = 10'h038;
        mem[373] = 10'h050;
        mem[374] = 10'h2f1;
        mem[375] = 10'h00a;
        mem[376] = 10'h008;
        mem[377] = 10'h29e;
        mem[378] = 10'h29b;
        mem[379] = 10'h3f7;
        mem[380] = 10'h0a3;
        mem[381] = 10'h176;
        mem[382] = 10'h38d;
        mem[383] = 10'h0ce;
        mem[384] = 10'h2c7;
        mem[385] = 10'h0fd;
        mem[386] = 10'h252;
        mem[387] = 10'h314;
        mem[388] = 10'h142;
        mem[389] = 10'h282;
        mem[390] = 10'h30d;
        mem[391] = 10'h19b;
        mem[392] = 10'h02c;
        mem[393] = 10'h086;
        mem[394] = 10'h260;
        mem[395] = 10'h3b6;
        mem[396] = 10'h357;
        mem[397] = 10'h22b;
        mem[398] = 10'h11c;
        mem[399] = 10'h363;
        mem[400] = 10'h1ba;
        mem[401] = 10'h07f;
        mem[402] = 10'h303;
        mem[403] = 10'h3c5;
        mem[404] = 10'h17d;
        mem[405] = 10'h274;
        mem[406] = 10'h1ce;
        mem[407] = 10'h141;
        mem[408] = 10'h062;
        mem[409] = 10'h3a5;
        mem[410] = 10'h1ef;
        mem[411] = 10'h06e;
        mem[412] = 10'h2e2;
        mem[413] = 10'h2f9;
        mem[414] = 10'h1e8;
        mem[415] = 10'h37a;
        mem[416] = 10'h1b3;
        mem[417] = 10'h2e3;
        mem[418] = 10'h04f;
        mem[419] = 10'h38a;
        mem[420] = 10'h16a;
        mem[421] = 10'h214;
        mem[422] = 10'h3bc;
        mem[423] = 10'h02e;
        mem[424] = 10'h2de;
        mem[425] = 10'h1c1;
        mem[426] = 10'h0e5;
        mem[427] = 10'h10b;
        mem[428] = 10'h28d;
        mem[429] = 10'h021;
        mem[430] = 10'h3be;
        mem[431] = 10'h20f;
        mem[432] = 10'h1a4;
        mem[433] = 10'h0ab;
        mem[434] = 10'h0e4;
        mem[435] = 10'h0b7;
        mem[436] = 10'h182;
        mem[437] = 10'h360;
        mem[438] = 10'h379;
        mem[439] = 10'h0bf;
        mem[440] = 10'h0d4;
        mem[441] = 10'h140;
        mem[442] = 10'h1da;
        mem[443] = 10'h1be;
        mem[444] = 10'h22d;
        mem[445] = 10'h185;
        mem[446] = 10'h068;
        mem[447] = 10'h031;
        mem[448] = 10'h00f;
        mem[449] = 10'h201;
        mem[450] = 10'h21f;
        mem[451] = 10'h31d;
        mem[452] = 10'h351;
        mem[453] = 10'h122;
        mem[454] = 10'h2ca;
        mem[455] = 10'h311;
        mem[456] = 10'h30b;
        mem[457] = 10'h250;
        mem[458] = 10'h20d;
        mem[459] = 10'h059;
        mem[460] = 10'h29f;
        mem[461] = 10'h01a;
        mem[462] = 10'h343;
        mem[463] = 10'h237;
        mem[464] = 10'h2e9;
        mem[465] = 10'h230;
        mem[466] = 10'h032;
        mem[467] = 10'h00e;
        mem[468] = 10'h196;
        mem[469] = 10'h040;
        mem[470] = 10'h1fb;
        mem[471] = 10'h261;
        mem[472] = 10'h046;
        mem[473] = 10'h16e;
        mem[474] = 10'h27d;
        mem[475] = 10'h296;
        mem[476] = 10'h1d5;
        mem[477] = 10'h264;
        mem[478] = 10'h07b;
        mem[479] = 10'h2b2;
        mem[480] = 10'h3e7;
        mem[481] = 10'h395;
        mem[482] = 10'h145;
        mem[483] = 10'h337;
        mem[484] = 10'h3c0;
        mem[485] = 10'h1ab;
        mem[486] = 10'h10f;
        mem[487] = 10'h25f;
        mem[488] = 10'h006;
        mem[489] = 10'h2f5;
        mem[490] = 10'h227;
        mem[491] = 10'h37d;
        mem[492] = 10'h070;
        mem[493] = 10'h0ef;
        mem[494] = 10'h139;
        mem[495] = 10'h1b9;
        mem[496] = 10'h365;
        mem[497] = 10'h2ae;
        mem[498] = 10'h2d4;
        mem[499] = 10'h0d1;
        mem[500] = 10'h101;
        mem[501] = 10'h228;
        mem[502] = 10'h067;
        mem[503] = 10'h25e;
        mem[504] = 10'h190;
        mem[505] = 10'h318;
        mem[506] = 10'h215;
        mem[507] = 10'h37f;
        mem[508] = 10'h2cb;
        mem[509] = 10'h1fd;
        mem[510] = 10'h168;
        mem[511] = 10'h3fb;
        mem[512] = 10'h270;
        mem[513] = 10'h3ab;
        mem[514] = 10'h3ad;
        mem[515] = 10'h053;
        mem[516] = 10'h1e7;
        mem[517] = 10'h299;
        mem[518] = 10'h018;
        mem[519] = 10'h331;
        mem[520] = 10'h255;
        mem[521] = 10'h287;
        mem[522] = 10'h104;
        mem[523] = 10'h1a1;
        mem[524] = 10'h28c;
        mem[525] = 10'h39c;
        mem[526] = 10'h08b;
        mem[527] = 10'h36e;
        mem[528] = 10'h263;
        mem[529] = 10'h118;
        mem[530] = 10'h315;
        mem[531] = 10'h302;
        mem[532] = 10'h3a3;
        mem[533] = 10'h244;
        mem[534] = 10'h010;
        mem[535] = 10'h33b;
        mem[536] = 10'h109;
        mem[537] = 10'h390;
        mem[538] = 10'h2e6;
        mem[539] = 10'h3f0;
        mem[540] = 10'h3ba;
        mem[541] = 10'h3f8;
        mem[542] = 10'h16f;
        mem[543] = 10'h3b3;
        mem[544] = 10'h017;
        mem[545] = 10'h2af;
        mem[546] = 10'h047;
        mem[547] = 10'h127;
        mem[548] = 10'h36f;
        mem[549] = 10'h0a1;
        mem[550] = 10'h1d3;
        mem[551] = 10'h175;
        mem[552] = 10'h2bd;
        mem[553] = 10'h224;
        mem[554] = 10'h133;
        mem[555] = 10'h21c;
        mem[556] = 10'h3a2;
        mem[557] = 10'h3da;
        mem[558] = 10'h097;
        mem[559] = 10'h21d;
        mem[560] = 10'h2f4;
        mem[561] = 10'h0c4;
        mem[562] = 10'h019;
        mem[563] = 10'h3d6;
        mem[564] = 10'h0c3;
        mem[565] = 10'h181;
        mem[566] = 10'h14b;
        mem[567] = 10'h0f3;
        mem[568] = 10'h353;
        mem[569] = 10'h2a2;
        mem[570] = 10'h08c;
        mem[571] = 10'h358;
        mem[572] = 10'h126;
        mem[573] = 10'h1ac;
        mem[574] = 10'h125;
        mem[575] = 10'h1e0;
        mem[576] = 10'h35c;
        mem[577] = 10'h2ee;
        mem[578] = 10'h11d;
        mem[579] = 10'h216;
        mem[580] = 10'h3db;
        mem[581] = 10'h073;
        mem[582] = 10'h348;
        mem[583] = 10'h391;
        mem[584] = 10'h100;
        mem[585] = 10'h301;
        mem[586] = 10'h2b0;
        mem[587] = 10'h012;
        mem[588] = 10'h1ad;
        mem[589] = 10'h039;
        mem[590] = 10'h3df;
        mem[591] = 10'h2ec;
        mem[592] = 10'h246;
        mem[593] = 10'h38e;
        mem[594] = 10'h096;
        mem[595] = 10'h19e;
        mem[596] = 10'h13c;
        mem[597] = 10'h2fa;
        mem[598] = 10'h36d;
        mem[599] = 10'h089;
        mem[600] = 10'h31b;
        mem[601] = 10'h05e;
        mem[602] = 10'h0cb;
        mem[603] = 10'h2a3;
        mem[604] = 10'h009;
        mem[605] = 10'h0a9;
        mem[606] = 10'h174;
        mem[607] = 10'h1c6;
        mem[608] = 10'h3ca;
        mem[609] = 10'h0a2;
        mem[610] = 10'h055;
        mem[611] = 10'h15b;
        mem[612] = 10'h0c6;
        mem[613] = 10'h350;
        mem[614] = 10'h1dd;
        mem[615] = 10'h1b6;
        mem[616] = 10'h0dc;
        mem[617] = 10'h361;
        mem[618] = 10'h0f9;
        mem[619] = 10'h24a;
        mem[620] = 10'h2b6;
        mem[621] = 10'h198;
        mem[622] = 10'h1a2;
        mem[623] = 10'h28e;
        mem[624] = 10'h1b2;
        mem[625] = 10'h0b0;
        mem[626] = 10'h3f9;
        mem[627] = 10'h31e;
        mem[628] = 10'h0b2;
        mem[629] = 10'h09b;
        mem[630] = 10'h0ac;
        mem[631] = 10'h2bc;
        mem[632] = 10'h31a;
        mem[633] = 10'h165;
        mem[634] = 10'h2b1;
        mem[635] = 10'h2d0;
        mem[636] = 10'h218;
        mem[637] = 10'h18f;
        mem[638] = 10'h2cc;
        mem[639] = 10'h2b4;
        mem[640] = 10'h026;
        mem[641] = 10'h1c9;
        mem[642] = 10'h211;
        mem[643] = 10'h24d;
        mem[644] = 10'h0f1;
        mem[645] = 10'h3ea;
        mem[646] = 10'h2a5;
        mem[647] = 10'h3fe;
        mem[648] = 10'h14c;
        mem[649] = 10'h35a;
        mem[650] = 10'h1e4;
        mem[651] = 10'h329;
        mem[652] = 10'h0df;
        mem[653] = 10'h09c;
        mem[654] = 10'h0d9;
        mem[655] = 10'h290;
        mem[656] = 10'h1dc;
        mem[657] = 10'h344;
        mem[658] = 10'h20c;
        mem[659] = 10'h3c7;
        mem[660] = 10'h3d0;
        mem[661] = 10'h2e5;
        mem[662] = 10'h19c;
        mem[663] = 10'h332;
        mem[664] = 10'h084;
        mem[665] = 10'h03c;
        mem[666] = 10'h3aa;
        mem[667] = 10'h072;
        mem[668] = 10'h0f5;
        mem[669] = 10'h103;
        mem[670] = 10'h0cf;
        mem[671] = 10'h0b1;
        mem[672] = 10'h03f;
        mem[673] = 10'h1d7;
        mem[674] = 10'h3e0;
        mem[675] = 10'h369;
        mem[676] = 10'h131;
        mem[677] = 10'h054;
        mem[678] = 10'h12c;
        mem[679] = 10'h0c5;
        mem[680] = 10'h370;
        mem[681] = 10'h098;
        mem[682] = 10'h3a0;
        mem[683] = 10'h085;
        mem[684] = 10'h3d8;
        mem[685] = 10'h0ff;
        mem[686] = 10'h1fc;
        mem[687] = 10'h1c7;
        mem[688] = 10'h1cb;
        mem[689] = 10'h2d2;
        mem[690] = 10'h0aa;
        mem[691] = 10'h352;
        mem[692] = 10'h108;
        mem[693] = 10'h149;
        mem[694] = 10'h312;
        mem[695] = 10'h18d;
        mem[696] = 10'h03d;
        mem[697] = 10'h071;
        mem[698] = 10'h1cf;
        mem[699] = 10'h2f2;
        mem[700] = 10'h0bc;
        mem[701] = 10'h1aa;
        mem[702] = 10'h2cd;
        mem[703] = 10'h160;
        mem[704] = 10'h25b;
        mem[705] = 10'h08f;
        mem[706] = 10'h19f;
        mem[707] = 10'h324;
        mem[708] = 10'h06f;
        mem[709] = 10'h277;
        mem[710] = 10'h138;
        mem[711] = 10'h367;
        mem[712] = 10'h234;
        mem[713] = 10'h157;
        mem[714] = 10'h197;
        mem[715] = 10'h2b9;
        mem[716] = 10'h3f6;
        mem[717] = 10'h289;
        mem[718] = 10'h3bd;
        mem[719] = 10'h049;
        mem[720] = 10'h080;
        mem[721] = 10'h05d;
        mem[722] = 10'h25c;
        mem[723] = 10'h0b8;
        mem[724] = 10'h24b;
        mem[725] = 10'h001;
        mem[726] = 10'h3c9;
        mem[727] = 10'h148;
        mem[728] = 10'h2b5;
        mem[729] = 10'h117;
        mem[730] = 10'h345;
        mem[731] = 10'h114;
        mem[732] = 10'h383;
        mem[733] = 10'h374;
        mem[734] = 10'h189;
        mem[735] = 10'h240;
        mem[736] = 10'h04c;
        mem[737] = 10'h2c1;
        mem[738] = 10'h041;
        mem[739] = 10'h317;
        mem[740] = 10'h0dd;
        mem[741] = 10'h39b;
        mem[742] = 10'h3c8;
        mem[743] = 10'h0f0;
        mem[744] = 10'h0ea;
        mem[745] = 10'h2ac;
        mem[746] = 10'h36b;
        mem[747] = 10'h015;
        mem[748] = 10'h136;
        mem[749] = 10'h04a;
        mem[750] = 10'h1c0;
        mem[751] = 10'h34f;
        mem[752] = 10'h003;
        mem[753] = 10'h23f;
        mem[754] = 10'h375;
        mem[755] = 10'h26e;
        mem[756] = 10'h12b;
        mem[757] = 10'h368;
        mem[758] = 10'h110;
        mem[759] = 10'h235;
        mem[760] = 10'h37b;
        mem[761] = 10'h123;
        mem[762] = 10'h11a;
        mem[763] = 10'h0d2;
        mem[764] = 10'h34d;
        mem[765] = 10'h27b;
        mem[766] = 10'h2fe;
        mem[767] = 10'h10e;
        mem[768] = 10'h06a;
        mem[769] = 10'h248;
        mem[770] = 10'h0da;
        mem[771] = 10'h076;
        mem[772] = 10'h293;
        mem[773] = 10'h1b1;
        mem[774] = 10'h191;
        mem[775] = 10'h30e;
        mem[776] = 10'h281;
        mem[777] = 10'h132;
        mem[778] = 10'h294;
        mem[779] = 10'h328;
        mem[780] = 10'h298;
        mem[781] = 10'h354;
        mem[782] = 10'h15d;
        mem[783] = 10'h38b;
        mem[784] = 10'h153;
        mem[785] = 10'h232;
        mem[786] = 10'h397;
        mem[787] = 10'h0fe;
        mem[788] = 10'h30f;
        mem[789] = 10'h048;
        mem[790] = 10'h3c6;
        mem[791] = 10'h24f;
        mem[792] = 10'h254;
        mem[793] = 10'h356;
        mem[794] = 10'h166;
        mem[795] = 10'h399;
        mem[796] = 10'h0cd;
        mem[797] = 10'h1e3;
        mem[798] = 10'h31f;
        mem[799] = 10'h135;
        mem[800] = 10'h0d8;
        mem[801] = 10'h074;
        mem[802] = 10'h0e1;
        mem[803] = 10'h01d;
        mem[804] = 10'h0e7;
        mem[805] = 10'h2d7;
        mem[806] = 10'h238;
        mem[807] = 10'h39a;
        mem[808] = 10'h241;
        mem[809] = 10'h0e0;
        mem[810] = 10'h17e;
        mem[811] = 10'h029;
        mem[812] = 10'h3a8;
        mem[813] = 10'h3b8;
        mem[814] = 10'h2db;
        mem[815] = 10'h0f8;
        mem[816] = 10'h116;
        mem[817] = 10'h3c3;
        mem[818] = 10'h05a;
        mem[819] = 10'h151;
        mem[820] = 10'h323;
        mem[821] = 10'h378;
        mem[822] = 10'h17b;
        mem[823] = 10'h3d2;
        mem[824] = 10'h327;
        mem[825] = 10'h15e;
        mem[826] = 10'h2c6;
        mem[827] = 10'h1d8;
        mem[828] = 10'h276;
        mem[829] = 10'h2cf;
        mem[830] = 10'h245;
        mem[831] = 10'h35b;
        mem[832] = 10'h180;
        mem[833] = 10'h1e6;
        mem[834] = 10'h0b9;
        mem[835] = 10'h3e2;
        mem[836] = 10'h033;
        mem[837] = 10'h335;
        mem[838] = 10'h262;
        mem[839] = 10'h042;
        mem[840] = 10'h233;
        mem[841] = 10'h128;
        mem[842] = 10'h007;
        mem[843] = 10'h04b;
        mem[844] = 10'h0c9;
        mem[845] = 10'h338;
        mem[846] = 10'h2fc;
        mem[847] = 10'h3b5;
        mem[848] = 10'h1d0;
        mem[849] = 10'h1eb;
        mem[850] = 10'h0bb;
        mem[851] = 10'h321;
        mem[852] = 10'h193;
        mem[853] = 10'h2e1;
        mem[854] = 10'h200;
        mem[855] = 10'h1ed;
        mem[856] = 10'h0ca;
        mem[857] = 10'h169;
        mem[858] = 10'h1a3;
        mem[859] = 10'h102;
        mem[860] = 10'h000;
        mem[861] = 10'h119;
        mem[862] = 10'h1ae;
        mem[863] = 10'h1bc;
        mem[864] = 10'h00d;
        mem[865] = 10'h25a;
        mem[866] = 10'h09f;
        mem[867] = 10'h371;
        mem[868] = 10'h2ce;
        mem[869] = 10'h313;
        mem[870] = 10'h115;
        mem[871] = 10'h1f9;
        mem[872] = 10'h1af;
        mem[873] = 10'h12d;
        mem[874] = 10'h3ac;
        mem[875] = 10'h01c;
        mem[876] = 10'h051;
        mem[877] = 10'h280;
        mem[878] = 10'h08a;
        mem[879] = 10'h381;
        mem[880] = 10'h212;
        mem[881] = 10'h0d6;
        mem[882] = 10'h060;
        mem[883] = 10'h1f7;
        mem[884] = 10'h33c;
        mem[885] = 10'h3c1;
        mem[886] = 10'h2f0;
        mem[887] = 10'h0f7;
        mem[888] = 10'h1bb;
        mem[889] = 10'h02f;
        mem[890] = 10'h056;
        mem[891] = 10'h095;
        mem[892] = 10'h3ef;
        mem[893] = 10'h326;
        mem[894] = 10'h23a;
        mem[895] = 10'h31c;
        mem[896] = 10'h20b;
        mem[897] = 10'h37e;
        mem[898] = 10'h1c4;
        mem[899] = 10'h0c2;
        mem[900] = 10'h2f3;
        mem[901] = 10'h265;
        mem[902] = 10'h088;
        mem[903] = 10'h32d;
        mem[904] = 10'h202;
        mem[905] = 10'h075;
        mem[906] = 10'h16c;
        mem[907] = 10'h023;
        mem[908] = 10'h07e;
        mem[909] = 10'h2a0;
        mem[910] = 10'h39d;
        mem[911] = 10'h164;
        mem[912] = 10'h09e;
        mem[913] = 10'h079;
        mem[914] = 10'h2bb;
        mem[915] = 10'h23e;
        mem[916] = 10'h0b3;
        mem[917] = 10'h155;
        mem[918] = 10'h13e;
        mem[919] = 10'h3e1;
        mem[920] = 10'h219;
        mem[921] = 10'h2d5;
        mem[922] = 10'h203;
        mem[923] = 10'h306;
        mem[924] = 10'h22f;
        mem[925] = 10'h0ed;
        mem[926] = 10'h347;
        mem[927] = 10'h1b0;
        mem[928] = 10'h147;
        mem[929] = 10'h078;
        mem[930] = 10'h2f7;
        mem[931] = 10'h077;
        mem[932] = 10'h01b;
        mem[933] = 10'h111;
        mem[934] = 10'h3e4;
        mem[935] = 10'h107;
        mem[936] = 10'h09d;
        mem[937] = 10'h39e;
        mem[938] = 10'h333;
        mem[939] = 10'h3d1;
        mem[940] = 10'h2b8;
        mem[941] = 10'h0c8;
        mem[942] = 10'h11b;
        mem[943] = 10'h1c2;
        mem[944] = 10'h025;
        mem[945] = 10'h016;
        mem[946] = 10'h207;
        mem[947] = 10'h386;
        mem[948] = 10'h011;
        mem[949] = 10'h1b7;
        mem[950] = 10'h18e;
        mem[951] = 10'h06c;
        mem[952] = 10'h284;
        mem[953] = 10'h3c4;
        mem[954] = 10'h130;
        mem[955] = 10'h063;
        mem[956] = 10'h002;
        mem[957] = 10'h0f4;
        mem[958] = 10'h3a4;
        mem[959] = 10'h129;
        mem[960] = 10'h1f8;
        mem[961] = 10'h194;
        mem[962] = 10'h06b;
        mem[963] = 10'h316;
        mem[964] = 10'h29c;
        mem[965] = 10'h087;
        mem[966] = 10'h339;
        mem[967] = 10'h33e;
        mem[968] = 10'h309;
        mem[969] = 10'h14d;
        mem[970] = 10'h178;
        mem[971] = 10'h3e6;
        mem[972] = 10'h08e;
        mem[973] = 10'h199;
        mem[974] = 10'h32a;
        mem[975] = 10'h39f;
        mem[976] = 10'h1c5;
        mem[977] = 10'h02b;
        mem[978] = 10'h13d;
        mem[979] = 10'h34a;
        mem[980] = 10'h0fc;
        mem[981] = 10'h1bf;
        mem[982] = 10'h13a;
        mem[983] = 10'h2ed;
        mem[984] = 10'h34c;
        mem[985] = 10'h0d3;
        mem[986] = 10'h307;
        mem[987] = 10'h156;
        mem[988] = 10'h1d4;
        mem[989] = 10'h3d3;
        mem[990] = 10'h1f3;
        mem[991] = 10'h179;
        mem[992] = 10'h1ec;
        mem[993] = 10'h2a8;
        mem[994] = 10'h06d;
        mem[995] = 10'h13b;
        mem[996] = 10'h035;
        mem[997] = 10'h09a;
        mem[998] = 10'h2df;
        mem[999] = 10'h394;
        mem[1000] = 10'h0fa;
        mem[1001] = 10'h2a6;
        mem[1002] = 10'h3dc;
        mem[1003] = 10'h32e;
        mem[1004] = 10'h02d;
        mem[1005] = 10'h295;
        mem[1006] = 10'h170;
        mem[1007] = 10'h161;
        mem[1008] = 10'h364;
        mem[1009] = 10'h398;
        mem[1010] = 10'h069;
        mem[1011] = 10'h2c8;
        mem[1012] = 10'h3af;
        mem[1013] = 10'h251;
        mem[1014] = 10'h04e;
        mem[1015] = 10'h19a;
        mem[1016] = 10'h1a5;
        mem[1017] = 10'h0bd;
        mem[1018] = 10'h093;
        mem[1019] = 10'h3b2;
        mem[1020] = 10'h028;
        mem[1021] = 10'h058;
        mem[1022] = 10'h037;
        mem[1023] = 10'h2d1;
    end
endmodule

module odo_apply_sboxes(clk, in, out);
    input clk;
    input [639:0] in;
    output [639:0] out;
    odo_sbox_small0 sbox0inst(clk, in[5:0], out[5:0]);
    odo_sbox_small1 sbox1inst(clk, in[21:16], out[21:16]);
    odo_sbox_large0 sbox2inst(clk, in[15:6], in[31:22], out[15:6], out[31:22]);
    odo_sbox_small2 sbox3inst(clk, in[37:32], out[37:32]);
    odo_sbox_small3 sbox4inst(clk, in[53:48], out[53:48]);
    odo_sbox_large0 sbox5inst(clk, in[47:38], in[63:54], out[47:38], out[63:54]);
    odo_sbox_small4 sbox6inst(clk, in[69:64], out[69:64]);
    odo_sbox_small5 sbox7inst(clk, in[85:80], out[85:80]);
    odo_sbox_large1 sbox8inst(clk, in[79:70], in[95:86], out[79:70], out[95:86]);
    odo_sbox_small6 sbox9inst(clk, in[101:96], out[101:96]);
    odo_sbox_small7 sbox10inst(clk, in[117:112], out[117:112]);
    odo_sbox_large1 sbox11inst(clk, in[111:102], in[127:118], out[111:102], out[127:118]);
    odo_sbox_small8 sbox12inst(clk, in[133:128], out[133:128]);
    odo_sbox_small9 sbox13inst(clk, in[149:144], out[149:144]);
    odo_sbox_large2 sbox14inst(clk, in[143:134], in[159:150], out[143:134], out[159:150]);
    odo_sbox_small10 sbox15inst(clk, in[165:160], out[165:160]);
    odo_sbox_small11 sbox16inst(clk, in[181:176], out[181:176]);
    odo_sbox_large2 sbox17inst(clk, in[175:166], in[191:182], out[175:166], out[191:182]);
    odo_sbox_small12 sbox18inst(clk, in[197:192], out[197:192]);
    odo_sbox_small13 sbox19inst(clk, in[213:208], out[213:208]);
    odo_sbox_large3 sbox20inst(clk, in[207:198], in[223:214], out[207:198], out[223:214]);
    odo_sbox_small14 sbox21inst(clk, in[229:224], out[229:224]);
    odo_sbox_small15 sbox22inst(clk, in[245:240], out[245:240]);
    odo_sbox_large3 sbox23inst(clk, in[239:230], in[255:246], out[239:230], out[255:246]);
    odo_sbox_small16 sbox24inst(clk, in[261:256], out[261:256]);
    odo_sbox_small17 sbox25inst(clk, in[277:272], out[277:272]);
    odo_sbox_large4 sbox26inst(clk, in[271:262], in[287:278], out[271:262], out[287:278]);
    odo_sbox_small18 sbox27inst(clk, in[293:288], out[293:288]);
    odo_sbox_small19 sbox28inst(clk, in[309:304], out[309:304]);
    odo_sbox_large4 sbox29inst(clk, in[303:294], in[319:310], out[303:294], out[319:310]);
    odo_sbox_small20 sbox30inst(clk, in[325:320], out[325:320]);
    odo_sbox_small21 sbox31inst(clk, in[341:336], out[341:336]);
    odo_sbox_large5 sbox32inst(clk, in[335:326], in[351:342], out[335:326], out[351:342]);
    odo_sbox_small22 sbox33inst(clk, in[357:352], out[357:352]);
    odo_sbox_small23 sbox34inst(clk, in[373:368], out[373:368]);
    odo_sbox_large5 sbox35inst(clk, in[367:358], in[383:374], out[367:358], out[383:374]);
    odo_sbox_small24 sbox36inst(clk, in[389:384], out[389:384]);
    odo_sbox_small25 sbox37inst(clk, in[405:400], out[405:400]);
    odo_sbox_large6 sbox38inst(clk, in[399:390], in[415:406], out[399:390], out[415:406]);
    odo_sbox_small26 sbox39inst(clk, in[421:416], out[421:416]);
    odo_sbox_small27 sbox40inst(clk, in[437:432], out[437:432]);
    odo_sbox_large6 sbox41inst(clk, in[431:422], in[447:438], out[431:422], out[447:438]);
    odo_sbox_small28 sbox42inst(clk, in[453:448], out[453:448]);
    odo_sbox_small29 sbox43inst(clk, in[469:464], out[469:464]);
    odo_sbox_large7 sbox44inst(clk, in[463:454], in[479:470], out[463:454], out[479:470]);
    odo_sbox_small30 sbox45inst(clk, in[485:480], out[485:480]);
    odo_sbox_small31 sbox46inst(clk, in[501:496], out[501:496]);
    odo_sbox_large7 sbox47inst(clk, in[495:486], in[511:502], out[495:486], out[511:502]);
    odo_sbox_small32 sbox48inst(clk, in[517:512], out[517:512]);
    odo_sbox_small33 sbox49inst(clk, in[533:528], out[533:528]);
    odo_sbox_large8 sbox50inst(clk, in[527:518], in[543:534], out[527:518], out[543:534]);
    odo_sbox_small34 sbox51inst(clk, in[549:544], out[549:544]);
    odo_sbox_small35 sbox52inst(clk, in[565:560], out[565:560]);
    odo_sbox_large8 sbox53inst(clk, in[559:550], in[575:566], out[559:550], out[575:566]);
    odo_sbox_small36 sbox54inst(clk, in[581:576], out[581:576]);
    odo_sbox_small37 sbox55inst(clk, in[597:592], out[597:592]);
    odo_sbox_large9 sbox56inst(clk, in[591:582], in[607:598], out[591:582], out[607:598]);
    odo_sbox_small38 sbox57inst(clk, in[613:608], out[613:608]);
    odo_sbox_small39 sbox58inst(clk, in[629:624], out[629:624]);
    odo_sbox_large9 sbox59inst(clk, in[623:614], in[639:630], out[623:614], out[639:630]);
endmodule

module odo_apply_pbox0(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[610] = in[0];
    assign out[532] = in[1];
    assign out[583] = in[2];
    assign out[307] = in[3];
    assign out[37] = in[4];
    assign out[146] = in[5];
    assign out[374] = in[6];
    assign out[311] = in[7];
    assign out[6] = in[8];
    assign out[313] = in[9];
    assign out[133] = in[10];
    assign out[315] = in[11];
    assign out[50] = in[12];
    assign out[16] = in[13];
    assign out[560] = in[14];
    assign out[490] = in[15];
    assign out[389] = in[16];
    assign out[209] = in[17];
    assign out[38] = in[18];
    assign out[241] = in[19];
    assign out[200] = in[20];
    assign out[123] = in[21];
    assign out[150] = in[22];
    assign out[56] = in[23];
    assign out[466] = in[24];
    assign out[75] = in[25];
    assign out[201] = in[26];
    assign out[25] = in[27];
    assign out[250] = in[28];
    assign out[575] = in[29];
    assign out[576] = in[30];
    assign out[189] = in[31];
    assign out[474] = in[32];
    assign out[149] = in[33];
    assign out[338] = in[34];
    assign out[477] = in[35];
    assign out[276] = in[36];
    assign out[462] = in[37];
    assign out[12] = in[38];
    assign out[284] = in[39];
    assign out[494] = in[40];
    assign out[350] = in[41];
    assign out[136] = in[42];
    assign out[589] = in[43];
    assign out[469] = in[44];
    assign out[264] = in[45];
    assign out[96] = in[46];
    assign out[163] = in[47];
    assign out[240] = in[48];
    assign out[371] = in[49];
    assign out[117] = in[50];
    assign out[231] = in[51];
    assign out[413] = in[52];
    assign out[634] = in[53];
    assign out[121] = in[54];
    assign out[105] = in[55];
    assign out[59] = in[56];
    assign out[379] = in[57];
    assign out[380] = in[58];
    assign out[15] = in[59];
    assign out[122] = in[60];
    assign out[472] = in[61];
    assign out[562] = in[62];
    assign out[424] = in[63];
    assign out[454] = in[64];
    assign out[21] = in[65];
    assign out[566] = in[66];
    assign out[428] = in[67];
    assign out[521] = in[68];
    assign out[387] = in[69];
    assign out[353] = in[70];
    assign out[194] = in[71];
    assign out[183] = in[72];
    assign out[111] = in[73];
    assign out[254] = in[74];
    assign out[134] = in[75];
    assign out[622] = in[76];
    assign out[386] = in[77];
    assign out[578] = in[78];
    assign out[324] = in[79];
    assign out[78] = in[80];
    assign out[275] = in[81];
    assign out[549] = in[82];
    assign out[147] = in[83];
    assign out[242] = in[84];
    assign out[552] = in[85];
    assign out[72] = in[86];
    assign out[139] = in[87];
    assign out[435] = in[88];
    assign out[282] = in[89];
    assign out[526] = in[90];
    assign out[637] = in[91];
    assign out[286] = in[92];
    assign out[419] = in[93];
    assign out[235] = in[94];
    assign out[485] = in[95];
    assign out[94] = in[96];
    assign out[156] = in[97];
    assign out[162] = in[98];
    assign out[425] = in[99];
    assign out[358] = in[100];
    assign out[11] = in[101];
    assign out[213] = in[102];
    assign out[42] = in[103];
    assign out[422] = in[104];
    assign out[169] = in[105];
    assign out[165] = in[106];
    assign out[300] = in[107];
    assign out[417] = in[108];
    assign out[83] = in[109];
    assign out[108] = in[110];
    assign out[501] = in[111];
    assign out[34] = in[112];
    assign out[613] = in[113];
    assign out[308] = in[114];
    assign out[412] = in[115];
    assign out[102] = in[116];
    assign out[233] = in[117];
    assign out[294] = in[118];
    assign out[416] = in[119];
    assign out[301] = in[120];
    assign out[557] = in[121];
    assign out[341] = in[122];
    assign out[512] = in[123];
    assign out[318] = in[124];
    assign out[507] = in[125];
    assign out[499] = in[126];
    assign out[101] = in[127];
    assign out[317] = in[128];
    assign out[372] = in[129];
    assign out[625] = in[130];
    assign out[443] = in[131];
    assign out[22] = in[132];
    assign out[628] = in[133];
    assign out[269] = in[134];
    assign out[89] = in[135];
    assign out[261] = in[136];
    assign out[548] = in[137];
    assign out[381] = in[138];
    assign out[600] = in[139];
    assign out[497] = in[140];
    assign out[544] = in[141];
    assign out[603] = in[142];
    assign out[500] = in[143];
    assign out[385] = in[144];
    assign out[450] = in[145];
    assign out[306] = in[146];
    assign out[76] = in[147];
    assign out[373] = in[148];
    assign out[558] = in[149];
    assign out[391] = in[150];
    assign out[266] = in[151];
    assign out[142] = in[152];
    assign out[550] = in[153];
    assign out[289] = in[154];
    assign out[630] = in[155];
    assign out[636] = in[156];
    assign out[62] = in[157];
    assign out[283] = in[158];
    assign out[607] = in[159];
    assign out[320] = in[160];
    assign out[503] = in[161];
    assign out[465] = in[162];
    assign out[47] = in[163];
    assign out[263] = in[164];
    assign out[406] = in[165];
    assign out[120] = in[166];
    assign out[112] = in[167];
    assign out[328] = in[168];
    assign out[329] = in[169];
    assign out[567] = in[170];
    assign out[267] = in[171];
    assign out[335] = in[172];
    assign out[246] = in[173];
    assign out[486] = in[174];
    assign out[181] = in[175];
    assign out[337] = in[176];
    assign out[509] = in[177];
    assign out[357] = in[178];
    assign out[518] = in[179];
    assign out[473] = in[180];
    assign out[190] = in[181];
    assign out[8] = in[182];
    assign out[382] = in[183];
    assign out[68] = in[184];
    assign out[255] = in[185];
    assign out[91] = in[186];
    assign out[455] = in[187];
    assign out[533] = in[188];
    assign out[536] = in[189];
    assign out[606] = in[190];
    assign out[32] = in[191];
    assign out[73] = in[192];
    assign out[64] = in[193];
    assign out[427] = in[194];
    assign out[214] = in[195];
    assign out[77] = in[196];
    assign out[268] = in[197];
    assign out[252] = in[198];
    assign out[360] = in[199];
    assign out[81] = in[200];
    assign out[298] = in[201];
    assign out[157] = in[202];
    assign out[481] = in[203];
    assign out[187] = in[204];
    assign out[110] = in[205];
    assign out[7] = in[206];
    assign out[48] = in[207];
    assign out[28] = in[208];
    assign out[344] = in[209];
    assign out[129] = in[210];
    assign out[166] = in[211];
    assign out[623] = in[212];
    assign out[196] = in[213];
    assign out[375] = in[214];
    assign out[160] = in[215];
    assign out[23] = in[216];
    assign out[238] = in[217];
    assign out[144] = in[218];
    assign out[448] = in[219];
    assign out[395] = in[220];
    assign out[554] = in[221];
    assign out[167] = in[222];
    assign out[40] = in[223];
    assign out[408] = in[224];
    assign out[170] = in[225];
    assign out[52] = in[226];
    assign out[611] = in[227];
    assign out[247] = in[228];
    assign out[184] = in[229];
    assign out[498] = in[230];
    assign out[615] = in[231];
    assign out[158] = in[232];
    assign out[585] = in[233];
    assign out[349] = in[234];
    assign out[270] = in[235];
    assign out[191] = in[236];
    assign out[520] = in[237];
    assign out[55] = in[238];
    assign out[274] = in[239];
    assign out[523] = in[240];
    assign out[198] = in[241];
    assign out[197] = in[242];
    assign out[491] = in[243];
    assign out[547] = in[244];
    assign out[528] = in[245];
    assign out[278] = in[246];
    assign out[599] = in[247];
    assign out[496] = in[248];
    assign out[601] = in[249];
    assign out[519] = in[250];
    assign out[302] = in[251];
    assign out[402] = in[252];
    assign out[60] = in[253];
    assign out[132] = in[254];
    assign out[459] = in[255];
    assign out[4] = in[256];
    assign out[69] = in[257];
    assign out[393] = in[258];
    assign out[423] = in[259];
    assign out[495] = in[260];
    assign out[45] = in[261];
    assign out[171] = in[262];
    assign out[343] = in[263];
    assign out[492] = in[264];
    assign out[620] = in[265];
    assign out[540] = in[266];
    assign out[363] = in[267];
    assign out[332] = in[268];
    assign out[41] = in[269];
    assign out[561] = in[270];
    assign out[249] = in[271];
    assign out[367] = in[272];
    assign out[394] = in[273];
    assign out[164] = in[274];
    assign out[116] = in[275];
    assign out[447] = in[276];
    assign out[483] = in[277];
    assign out[310] = in[278];
    assign out[130] = in[279];
    assign out[571] = in[280];
    assign out[281] = in[281];
    assign out[346] = in[282];
    assign out[128] = in[283];
    assign out[206] = in[284];
    assign out[135] = in[285];
    assign out[591] = in[286];
    assign out[280] = in[287];
    assign out[138] = in[288];
    assign out[243] = in[289];
    assign out[543] = in[290];
    assign out[323] = in[291];
    assign out[348] = in[292];
    assign out[464] = in[293];
    assign out[152] = in[294];
    assign out[145] = in[295];
    assign out[570] = in[296];
    assign out[432] = in[297];
    assign out[546] = in[298];
    assign out[399] = in[299];
    assign out[293] = in[300];
    assign out[151] = in[301];
    assign out[437] = in[302];
    assign out[30] = in[303];
    assign out[218] = in[304];
    assign out[476] = in[305];
    assign out[19] = in[306];
    assign out[605] = in[307];
    assign out[205] = in[308];
    assign out[154] = in[309];
    assign out[277] = in[310];
    assign out[95] = in[311];
    assign out[390] = in[312];
    assign out[384] = in[313];
    assign out[612] = in[314];
    assign out[106] = in[315];
    assign out[36] = in[316];
    assign out[155] = in[317];
    assign out[418] = in[318];
    assign out[504] = in[319];
    assign out[178] = in[320];
    assign out[257] = in[321];
    assign out[322] = in[322];
    assign out[245] = in[323];
    assign out[598] = in[324];
    assign out[9] = in[325];
    assign out[426] = in[326];
    assign out[618] = in[327];
    assign out[256] = in[328];
    assign out[265] = in[329];
    assign out[239] = in[330];
    assign out[58] = in[331];
    assign out[299] = in[332];
    assign out[230] = in[333];
    assign out[505] = in[334];
    assign out[626] = in[335];
    assign out[186] = in[336];
    assign out[109] = in[337];
    assign out[290] = in[338];
    assign out[488] = in[339];
    assign out[631] = in[340];
    assign out[551] = in[341];
    assign out[342] = in[342];
    assign out[279] = in[343];
    assign out[0] = in[344];
    assign out[619] = in[345];
    assign out[179] = in[346];
    assign out[124] = in[347];
    assign out[639] = in[348];
    assign out[316] = in[349];
    assign out[584] = in[350];
    assign out[14] = in[351];
    assign out[487] = in[352];
    assign out[587] = in[353];
    assign out[126] = in[354];
    assign out[63] = in[355];
    assign out[5] = in[356];
    assign out[414] = in[357];
    assign out[493] = in[358];
    assign out[43] = in[359];
    assign out[312] = in[360];
    assign out[297] = in[361];
    assign out[398] = in[362];
    assign out[616] = in[363];
    assign out[292] = in[364];
    assign out[542] = in[365];
    assign out[10] = in[366];
    assign out[530] = in[367];
    assign out[545] = in[368];
    assign out[18] = in[369];
    assign out[258] = in[370];
    assign out[119] = in[371];
    assign out[35] = in[372];
    assign out[57] = in[373];
    assign out[82] = in[374];
    assign out[137] = in[375];
    assign out[20] = in[376];
    assign out[104] = in[377];
    assign out[216] = in[378];
    assign out[436] = in[379];
    assign out[480] = in[380];
    assign out[175] = in[381];
    assign out[334] = in[382];
    assign out[228] = in[383];
    assign out[340] = in[384];
    assign out[527] = in[385];
    assign out[207] = in[386];
    assign out[79] = in[387];
    assign out[522] = in[388];
    assign out[211] = in[389];
    assign out[354] = in[390];
    assign out[273] = in[391];
    assign out[118] = in[392];
    assign out[143] = in[393];
    assign out[345] = in[394];
    assign out[525] = in[395];
    assign out[579] = in[396];
    assign out[29] = in[397];
    assign out[215] = in[398];
    assign out[597] = in[399];
    assign out[330] = in[400];
    assign out[515] = in[401];
    assign out[159] = in[402];
    assign out[1] = in[403];
    assign out[225] = in[404];
    assign out[535] = in[405];
    assign out[430] = in[406];
    assign out[452] = in[407];
    assign out[80] = in[408];
    assign out[539] = in[409];
    assign out[224] = in[410];
    assign out[362] = in[411];
    assign out[226] = in[412];
    assign out[88] = in[413];
    assign out[46] = in[414];
    assign out[90] = in[415];
    assign out[24] = in[416];
    assign out[559] = in[417];
    assign out[114] = in[418];
    assign out[319] = in[419];
    assign out[608] = in[420];
    assign out[221] = in[421];
    assign out[236] = in[422];
    assign out[638] = in[423];
    assign out[444] = in[424];
    assign out[555] = in[425];
    assign out[98] = in[426];
    assign out[309] = in[427];
    assign out[409] = in[428];
    assign out[449] = in[429];
    assign out[624] = in[430];
    assign out[451] = in[431];
    assign out[260] = in[432];
    assign out[441] = in[433];
    assign out[251] = in[434];
    assign out[33] = in[435];
    assign out[336] = in[436];
    assign out[383] = in[437];
    assign out[174] = in[438];
    assign out[321] = in[439];
    assign out[582] = in[440];
    assign out[333] = in[441];
    assign out[457] = in[442];
    assign out[467] = in[443];
    assign out[232] = in[444];
    assign out[53] = in[445];
    assign out[204] = in[446];
    assign out[471] = in[447];
    assign out[271] = in[448];
    assign out[173] = in[449];
    assign out[203] = in[450];
    assign out[44] = in[451];
    assign out[403] = in[452];
    assign out[604] = in[453];
    assign out[405] = in[454];
    assign out[2] = in[455];
    assign out[407] = in[456];
    assign out[339] = in[457];
    assign out[577] = in[458];
    assign out[593] = in[459];
    assign out[484] = in[460];
    assign out[219] = in[461];
    assign out[596] = in[462];
    assign out[478] = in[463];
    assign out[364] = in[464];
    assign out[17] = in[465];
    assign out[202] = in[466];
    assign out[295] = in[467];
    assign out[592] = in[468];
    assign out[13] = in[469];
    assign out[227] = in[470];
    assign out[531] = in[471];
    assign out[538] = in[472];
    assign out[223] = in[473];
    assign out[361] = in[474];
    assign out[303] = in[475];
    assign out[212] = in[476];
    assign out[70] = in[477];
    assign out[556] = in[478];
    assign out[396] = in[479];
    assign out[27] = in[480];
    assign out[632] = in[481];
    assign out[442] = in[482];
    assign out[602] = in[483];
    assign out[234] = in[484];
    assign out[287] = in[485];
    assign out[244] = in[486];
    assign out[369] = in[487];
    assign out[148] = in[488];
    assign out[440] = in[489];
    assign out[568] = in[490];
    assign out[506] = in[491];
    assign out[103] = in[492];
    assign out[410] = in[493];
    assign out[502] = in[494];
    assign out[446] = in[495];
    assign out[388] = in[496];
    assign out[563] = in[497];
    assign out[326] = in[498];
    assign out[586] = in[499];
    assign out[93] = in[500];
    assign out[445] = in[501];
    assign out[31] = in[502];
    assign out[463] = in[503];
    assign out[370] = in[504];
    assign out[259] = in[505];
    assign out[529] = in[506];
    assign out[100] = in[507];
    assign out[180] = in[508];
    assign out[327] = in[509];
    assign out[39] = in[510];
    assign out[140] = in[511];
    assign out[172] = in[512];
    assign out[581] = in[513];
    assign out[176] = in[514];
    assign out[415] = in[515];
    assign out[107] = in[516];
    assign out[633] = in[517];
    assign out[400] = in[518];
    assign out[125] = in[519];
    assign out[524] = in[520];
    assign out[352] = in[521];
    assign out[325] = in[522];
    assign out[188] = in[523];
    assign out[331] = in[524];
    assign out[513] = in[525];
    assign out[49] = in[526];
    assign out[253] = in[527];
    assign out[580] = in[528];
    assign out[569] = in[529];
    assign out[131] = in[530];
    assign out[516] = in[531];
    assign out[489] = in[532];
    assign out[185] = in[533];
    assign out[574] = in[534];
    assign out[517] = in[535];
    assign out[482] = in[536];
    assign out[304] = in[537];
    assign out[537] = in[538];
    assign out[74] = in[539];
    assign out[3] = in[540];
    assign out[65] = in[541];
    assign out[588] = in[542];
    assign out[141] = in[543];
    assign out[347] = in[544];
    assign out[288] = in[545];
    assign out[195] = in[546];
    assign out[272] = in[547];
    assign out[420] = in[548];
    assign out[617] = in[549];
    assign out[397] = in[550];
    assign out[291] = in[551];
    assign out[534] = in[552];
    assign out[356] = in[553];
    assign out[511] = in[554];
    assign out[431] = in[555];
    assign out[392] = in[556];
    assign out[217] = in[557];
    assign out[621] = in[558];
    assign out[86] = in[559];
    assign out[222] = in[560];
    assign out[84] = in[561];
    assign out[97] = in[562];
    assign out[161] = in[563];
    assign out[475] = in[564];
    assign out[401] = in[565];
    assign out[438] = in[566];
    assign out[229] = in[567];
    assign out[177] = in[568];
    assign out[609] = in[569];
    assign out[510] = in[570];
    assign out[553] = in[571];
    assign out[168] = in[572];
    assign out[351] = in[573];
    assign out[378] = in[574];
    assign out[314] = in[575];
    assign out[564] = in[576];
    assign out[453] = in[577];
    assign out[113] = in[578];
    assign out[461] = in[579];
    assign out[629] = in[580];
    assign out[439] = in[581];
    assign out[411] = in[582];
    assign out[565] = in[583];
    assign out[572] = in[584];
    assign out[237] = in[585];
    assign out[479] = in[586];
    assign out[627] = in[587];
    assign out[115] = in[588];
    assign out[67] = in[589];
    assign out[514] = in[590];
    assign out[192] = in[591];
    assign out[51] = in[592];
    assign out[71] = in[593];
    assign out[54] = in[594];
    assign out[635] = in[595];
    assign out[248] = in[596];
    assign out[193] = in[597];
    assign out[285] = in[598];
    assign out[208] = in[599];
    assign out[458] = in[600];
    assign out[61] = in[601];
    assign out[590] = in[602];
    assign out[127] = in[603];
    assign out[433] = in[604];
    assign out[434] = in[605];
    assign out[541] = in[606];
    assign out[66] = in[607];
    assign out[153] = in[608];
    assign out[421] = in[609];
    assign out[404] = in[610];
    assign out[199] = in[611];
    assign out[470] = in[612];
    assign out[595] = in[613];
    assign out[365] = in[614];
    assign out[366] = in[615];
    assign out[87] = in[616];
    assign out[368] = in[617];
    assign out[594] = in[618];
    assign out[220] = in[619];
    assign out[359] = in[620];
    assign out[429] = in[621];
    assign out[210] = in[622];
    assign out[262] = in[623];
    assign out[460] = in[624];
    assign out[85] = in[625];
    assign out[508] = in[626];
    assign out[456] = in[627];
    assign out[99] = in[628];
    assign out[305] = in[629];
    assign out[355] = in[630];
    assign out[26] = in[631];
    assign out[614] = in[632];
    assign out[92] = in[633];
    assign out[377] = in[634];
    assign out[296] = in[635];
    assign out[376] = in[636];
    assign out[182] = in[637];
    assign out[573] = in[638];
    assign out[468] = in[639];
endmodule

module odo_apply_pbox1(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[48] = in[0];
    assign out[613] = in[1];
    assign out[130] = in[2];
    assign out[242] = in[3];
    assign out[71] = in[4];
    assign out[157] = in[5];
    assign out[73] = in[6];
    assign out[294] = in[7];
    assign out[571] = in[8];
    assign out[419] = in[9];
    assign out[41] = in[10];
    assign out[588] = in[11];
    assign out[422] = in[12];
    assign out[125] = in[13];
    assign out[304] = in[14];
    assign out[143] = in[15];
    assign out[256] = in[16];
    assign out[536] = in[17];
    assign out[308] = in[18];
    assign out[371] = in[19];
    assign out[583] = in[20];
    assign out[633] = in[21];
    assign out[38] = in[22];
    assign out[151] = in[23];
    assign out[403] = in[24];
    assign out[545] = in[25];
    assign out[539] = in[26];
    assign out[43] = in[27];
    assign out[268] = in[28];
    assign out[238] = in[29];
    assign out[381] = in[30];
    assign out[280] = in[31];
    assign out[411] = in[32];
    assign out[546] = in[33];
    assign out[518] = in[34];
    assign out[115] = in[35];
    assign out[319] = in[36];
    assign out[557] = in[37];
    assign out[586] = in[38];
    assign out[385] = in[39];
    assign out[344] = in[40];
    assign out[561] = in[41];
    assign out[438] = in[42];
    assign out[203] = in[43];
    assign out[543] = in[44];
    assign out[156] = in[45];
    assign out[72] = in[46];
    assign out[334] = in[47];
    assign out[113] = in[48];
    assign out[50] = in[49];
    assign out[547] = in[50];
    assign out[461] = in[51];
    assign out[197] = in[52];
    assign out[302] = in[53];
    assign out[450] = in[54];
    assign out[16] = in[55];
    assign out[501] = in[56];
    assign out[570] = in[57];
    assign out[233] = in[58];
    assign out[579] = in[59];
    assign out[220] = in[60];
    assign out[638] = in[61];
    assign out[150] = in[62];
    assign out[350] = in[63];
    assign out[377] = in[64];
    assign out[288] = in[65];
    assign out[429] = in[66];
    assign out[195] = in[67];
    assign out[228] = in[68];
    assign out[401] = in[69];
    assign out[433] = in[70];
    assign out[152] = in[71];
    assign out[585] = in[72];
    assign out[248] = in[73];
    assign out[357] = in[74];
    assign out[260] = in[75];
    assign out[502] = in[76];
    assign out[596] = in[77];
    assign out[104] = in[78];
    assign out[534] = in[79];
    assign out[47] = in[80];
    assign out[321] = in[81];
    assign out[445] = in[82];
    assign out[86] = in[83];
    assign out[229] = in[84];
    assign out[584] = in[85];
    assign out[496] = in[86];
    assign out[606] = in[87];
    assign out[49] = in[88];
    assign out[602] = in[89];
    assign out[339] = in[90];
    assign out[310] = in[91];
    assign out[390] = in[92];
    assign out[392] = in[93];
    assign out[182] = in[94];
    assign out[505] = in[95];
    assign out[616] = in[96];
    assign out[532] = in[97];
    assign out[258] = in[98];
    assign out[251] = in[99];
    assign out[67] = in[100];
    assign out[189] = in[101];
    assign out[262] = in[102];
    assign out[465] = in[103];
    assign out[215] = in[104];
    assign out[281] = in[105];
    assign out[452] = in[106];
    assign out[252] = in[107];
    assign out[487] = in[108];
    assign out[173] = in[109];
    assign out[427] = in[110];
    assign out[239] = in[111];
    assign out[74] = in[112];
    assign out[569] = in[113];
    assign out[146] = in[114];
    assign out[162] = in[115];
    assign out[635] = in[116];
    assign out[245] = in[117];
    assign out[499] = in[118];
    assign out[103] = in[119];
    assign out[512] = in[120];
    assign out[217] = in[121];
    assign out[341] = in[122];
    assign out[60] = in[123];
    assign out[141] = in[124];
    assign out[285] = in[125];
    assign out[237] = in[126];
    assign out[2] = in[127];
    assign out[589] = in[128];
    assign out[359] = in[129];
    assign out[423] = in[130];
    assign out[116] = in[131];
    assign out[553] = in[132];
    assign out[98] = in[133];
    assign out[485] = in[134];
    assign out[180] = in[135];
    assign out[188] = in[136];
    assign out[391] = in[137];
    assign out[59] = in[138];
    assign out[420] = in[139];
    assign out[421] = in[140];
    assign out[241] = in[141];
    assign out[526] = in[142];
    assign out[444] = in[143];
    assign out[270] = in[144];
    assign out[336] = in[145];
    assign out[607] = in[146];
    assign out[626] = in[147];
    assign out[378] = in[148];
    assign out[573] = in[149];
    assign out[7] = in[150];
    assign out[81] = in[151];
    assign out[484] = in[152];
    assign out[550] = in[153];
    assign out[57] = in[154];
    assign out[348] = in[155];
    assign out[347] = in[156];
    assign out[517] = in[157];
    assign out[503] = in[158];
    assign out[413] = in[159];
    assign out[196] = in[160];
    assign out[565] = in[161];
    assign out[328] = in[162];
    assign out[0] = in[163];
    assign out[85] = in[164];
    assign out[291] = in[165];
    assign out[332] = in[166];
    assign out[123] = in[167];
    assign out[297] = in[168];
    assign out[6] = in[169];
    assign out[527] = in[170];
    assign out[361] = in[171];
    assign out[224] = in[172];
    assign out[364] = in[173];
    assign out[31] = in[174];
    assign out[493] = in[175];
    assign out[399] = in[176];
    assign out[581] = in[177];
    assign out[99] = in[178];
    assign out[447] = in[179];
    assign out[37] = in[180];
    assign out[449] = in[181];
    assign out[19] = in[182];
    assign out[349] = in[183];
    assign out[541] = in[184];
    assign out[508] = in[185];
    assign out[601] = in[186];
    assign out[289] = in[187];
    assign out[27] = in[188];
    assign out[476] = in[189];
    assign out[605] = in[190];
    assign out[428] = in[191];
    assign out[396] = in[192];
    assign out[533] = in[193];
    assign out[166] = in[194];
    assign out[32] = in[195];
    assign out[489] = in[196];
    assign out[498] = in[197];
    assign out[530] = in[198];
    assign out[486] = in[199];
    assign out[201] = in[200];
    assign out[494] = in[201];
    assign out[174] = in[202];
    assign out[393] = in[203];
    assign out[240] = in[204];
    assign out[464] = in[205];
    assign out[271] = in[206];
    assign out[402] = in[207];
    assign out[568] = in[208];
    assign out[311] = in[209];
    assign out[511] = in[210];
    assign out[4] = in[211];
    assign out[435] = in[212];
    assign out[269] = in[213];
    assign out[598] = in[214];
    assign out[535] = in[215];
    assign out[119] = in[216];
    assign out[253] = in[217];
    assign out[578] = in[218];
    assign out[136] = in[219];
    assign out[340] = in[220];
    assign out[124] = in[221];
    assign out[88] = in[222];
    assign out[147] = in[223];
    assign out[483] = in[224];
    assign out[206] = in[225];
    assign out[480] = in[226];
    assign out[386] = in[227];
    assign out[120] = in[228];
    assign out[121] = in[229];
    assign out[138] = in[230];
    assign out[333] = in[231];
    assign out[132] = in[232];
    assign out[158] = in[233];
    assign out[463] = in[234];
    assign out[298] = in[235];
    assign out[29] = in[236];
    assign out[293] = in[237];
    assign out[226] = in[238];
    assign out[163] = in[239];
    assign out[15] = in[240];
    assign out[34] = in[241];
    assign out[395] = in[242];
    assign out[100] = in[243];
    assign out[537] = in[244];
    assign out[301] = in[245];
    assign out[266] = in[246];
    assign out[40] = in[247];
    assign out[23] = in[248];
    assign out[221] = in[249];
    assign out[222] = in[250];
    assign out[53] = in[251];
    assign out[379] = in[252];
    assign out[177] = in[253];
    assign out[477] = in[254];
    assign out[92] = in[255];
    assign out[212] = in[256];
    assign out[560] = in[257];
    assign out[322] = in[258];
    assign out[318] = in[259];
    assign out[231] = in[260];
    assign out[513] = in[261];
    assign out[10] = in[262];
    assign out[155] = in[263];
    assign out[83] = in[264];
    assign out[367] = in[265];
    assign out[360] = in[266];
    assign out[25] = in[267];
    assign out[425] = in[268];
    assign out[89] = in[269];
    assign out[637] = in[270];
    assign out[398] = in[271];
    assign out[243] = in[272];
    assign out[576] = in[273];
    assign out[94] = in[274];
    assign out[504] = in[275];
    assign out[168] = in[276];
    assign out[516] = in[277];
    assign out[636] = in[278];
    assign out[317] = in[279];
    assign out[548] = in[280];
    assign out[101] = in[281];
    assign out[416] = in[282];
    assign out[577] = in[283];
    assign out[441] = in[284];
    assign out[442] = in[285];
    assign out[129] = in[286];
    assign out[179] = in[287];
    assign out[453] = in[288];
    assign out[45] = in[289];
    assign out[603] = in[290];
    assign out[295] = in[291];
    assign out[292] = in[292];
    assign out[625] = in[293];
    assign out[358] = in[294];
    assign out[114] = in[295];
    assign out[54] = in[296];
    assign out[440] = in[297];
    assign out[198] = in[298];
    assign out[106] = in[299];
    assign out[457] = in[300];
    assign out[137] = in[301];
    assign out[164] = in[302];
    assign out[58] = in[303];
    assign out[140] = in[304];
    assign out[133] = in[305];
    assign out[287] = in[306];
    assign out[345] = in[307];
    assign out[234] = in[308];
    assign out[509] = in[309];
    assign out[514] = in[310];
    assign out[329] = in[311];
    assign out[628] = in[312];
    assign out[205] = in[313];
    assign out[352] = in[314];
    assign out[118] = in[315];
    assign out[473] = in[316];
    assign out[209] = in[317];
    assign out[244] = in[318];
    assign out[126] = in[319];
    assign out[456] = in[320];
    assign out[384] = in[321];
    assign out[165] = in[322];
    assign out[185] = in[323];
    assign out[8] = in[324];
    assign out[9] = in[325];
    assign out[82] = in[326];
    assign out[66] = in[327];
    assign out[462] = in[328];
    assign out[191] = in[329];
    assign out[149] = in[330];
    assign out[580] = in[331];
    assign out[520] = in[332];
    assign out[351] = in[333];
    assign out[491] = in[334];
    assign out[587] = in[335];
    assign out[20] = in[336];
    assign out[574] = in[337];
    assign out[632] = in[338];
    assign out[466] = in[339];
    assign out[528] = in[340];
    assign out[307] = in[341];
    assign out[323] = in[342];
    assign out[343] = in[343];
    assign out[172] = in[344];
    assign out[408] = in[345];
    assign out[376] = in[346];
    assign out[183] = in[347];
    assign out[265] = in[348];
    assign out[192] = in[349];
    assign out[286] = in[350];
    assign out[194] = in[351];
    assign out[382] = in[352];
    assign out[44] = in[353];
    assign out[112] = in[354];
    assign out[559] = in[355];
    assign out[128] = in[356];
    assign out[523] = in[357];
    assign out[562] = in[358];
    assign out[460] = in[359];
    assign out[51] = in[360];
    assign out[600] = in[361];
    assign out[380] = in[362];
    assign out[400] = in[363];
    assign out[207] = in[364];
    assign out[538] = in[365];
    assign out[122] = in[366];
    assign out[61] = in[367];
    assign out[111] = in[368];
    assign out[406] = in[369];
    assign out[134] = in[370];
    assign out[169] = in[371];
    assign out[303] = in[372];
    assign out[388] = in[373];
    assign out[202] = in[374];
    assign out[211] = in[375];
    assign out[542] = in[376];
    assign out[213] = in[377];
    assign out[563] = in[378];
    assign out[609] = in[379];
    assign out[216] = in[380];
    assign out[620] = in[381];
    assign out[225] = in[382];
    assign out[219] = in[383];
    assign out[63] = in[384];
    assign out[64] = in[385];
    assign out[1] = in[386];
    assign out[624] = in[387];
    assign out[469] = in[388];
    assign out[608] = in[389];
    assign out[470] = in[390];
    assign out[610] = in[391];
    assign out[506] = in[392];
    assign out[443] = in[393];
    assign out[567] = in[394];
    assign out[273] = in[395];
    assign out[320] = in[396];
    assign out[12] = in[397];
    assign out[14] = in[398];
    assign out[277] = in[399];
    assign out[278] = in[400];
    assign out[482] = in[401];
    assign out[148] = in[402];
    assign out[621] = in[403];
    assign out[282] = in[404];
    assign out[558] = in[405];
    assign out[235] = in[406];
    assign out[267] = in[407];
    assign out[218] = in[408];
    assign out[159] = in[409];
    assign out[552] = in[410];
    assign out[492] = in[411];
    assign out[387] = in[412];
    assign out[199] = in[413];
    assign out[524] = in[414];
    assign out[454] = in[415];
    assign out[95] = in[416];
    assign out[96] = in[417];
    assign out[296] = in[418];
    assign out[78] = in[419];
    assign out[90] = in[420];
    assign out[160] = in[421];
    assign out[564] = in[422];
    assign out[108] = in[423];
    assign out[210] = in[424];
    assign out[599] = in[425];
    assign out[105] = in[426];
    assign out[368] = in[427];
    assign out[305] = in[428];
    assign out[109] = in[429];
    assign out[46] = in[430];
    assign out[372] = in[431];
    assign out[407] = in[432];
    assign out[375] = in[433];
    assign out[312] = in[434];
    assign out[181] = in[435];
    assign out[475] = in[436];
    assign out[315] = in[437];
    assign out[488] = in[438];
    assign out[612] = in[439];
    assign out[595] = in[440];
    assign out[56] = in[441];
    assign out[551] = in[442];
    assign out[144] = in[443];
    assign out[254] = in[444];
    assign out[284] = in[445];
    assign out[324] = in[446];
    assign out[556] = in[447];
    assign out[622] = in[448];
    assign out[131] = in[449];
    assign out[264] = in[450];
    assign out[110] = in[451];
    assign out[68] = in[452];
    assign out[69] = in[453];
    assign out[338] = in[454];
    assign out[544] = in[455];
    assign out[178] = in[456];
    assign out[566] = in[457];
    assign out[272] = in[458];
    assign out[65] = in[459];
    assign out[17] = in[460];
    assign out[275] = in[461];
    assign out[208] = in[462];
    assign out[572] = in[463];
    assign out[21] = in[464];
    assign out[417] = in[465];
    assign out[619] = in[466];
    assign out[24] = in[467];
    assign out[127] = in[468];
    assign out[283] = in[469];
    assign out[290] = in[470];
    assign out[236] = in[471];
    assign out[394] = in[472];
    assign out[615] = in[473];
    assign out[519] = in[474];
    assign out[26] = in[475];
    assign out[353] = in[476];
    assign out[630] = in[477];
    assign out[356] = in[478];
    assign out[36] = in[479];
    assign out[432] = in[480];
    assign out[467] = in[481];
    assign out[257] = in[482];
    assign out[405] = in[483];
    assign out[593] = in[484];
    assign out[91] = in[485];
    assign out[439] = in[486];
    assign out[84] = in[487];
    assign out[39] = in[488];
    assign out[631] = in[489];
    assign out[507] = in[490];
    assign out[582] = in[491];
    assign out[87] = in[492];
    assign out[232] = in[493];
    assign out[481] = in[494];
    assign out[153] = in[495];
    assign out[335] = in[496];
    assign out[374] = in[497];
    assign out[337] = in[498];
    assign out[313] = in[499];
    assign out[250] = in[500];
    assign out[389] = in[501];
    assign out[35] = in[502];
    assign out[342] = in[503];
    assign out[549] = in[504];
    assign out[255] = in[505];
    assign out[459] = in[506];
    assign out[418] = in[507];
    assign out[145] = in[508];
    assign out[369] = in[509];
    assign out[370] = in[510];
    assign out[525] = in[511];
    assign out[604] = in[512];
    assign out[184] = in[513];
    assign out[247] = in[514];
    assign out[437] = in[515];
    assign out[249] = in[516];
    assign out[597] = in[517];
    assign out[223] = in[518];
    assign out[79] = in[519];
    assign out[592] = in[520];
    assign out[529] = in[521];
    assign out[531] = in[522];
    assign out[227] = in[523];
    assign out[479] = in[524];
    assign out[230] = in[525];
    assign out[554] = in[526];
    assign out[555] = in[527];
    assign out[117] = in[528];
    assign out[451] = in[529];
    assign out[55] = in[530];
    assign out[500] = in[531];
    assign out[327] = in[532];
    assign out[204] = in[533];
    assign out[331] = in[534];
    assign out[62] = in[535];
    assign out[70] = in[536];
    assign out[629] = in[537];
    assign out[354] = in[538];
    assign out[397] = in[539];
    assign out[510] = in[540];
    assign out[75] = in[541];
    assign out[246] = in[542];
    assign out[623] = in[543];
    assign out[5] = in[544];
    assign out[436] = in[545];
    assign out[42] = in[546];
    assign out[187] = in[547];
    assign out[300] = in[548];
    assign out[154] = in[549];
    assign out[366] = in[550];
    assign out[346] = in[551];
    assign out[77] = in[552];
    assign out[80] = in[553];
    assign out[412] = in[554];
    assign out[627] = in[555];
    assign out[478] = in[556];
    assign out[448] = in[557];
    assign out[28] = in[558];
    assign out[93] = in[559];
    assign out[167] = in[560];
    assign out[276] = in[561];
    assign out[404] = in[562];
    assign out[170] = in[563];
    assign out[455] = in[564];
    assign out[142] = in[565];
    assign out[424] = in[566];
    assign out[409] = in[567];
    assign out[426] = in[568];
    assign out[410] = in[569];
    assign out[522] = in[570];
    assign out[316] = in[571];
    assign out[414] = in[572];
    assign out[495] = in[573];
    assign out[214] = in[574];
    assign out[97] = in[575];
    assign out[373] = in[576];
    assign out[468] = in[577];
    assign out[594] = in[578];
    assign out[11] = in[579];
    assign out[102] = in[580];
    assign out[314] = in[581];
    assign out[52] = in[582];
    assign out[190] = in[583];
    assign out[363] = in[584];
    assign out[107] = in[585];
    assign out[383] = in[586];
    assign out[306] = in[587];
    assign out[446] = in[588];
    assign out[614] = in[589];
    assign out[259] = in[590];
    assign out[279] = in[591];
    assign out[135] = in[592];
    assign out[618] = in[593];
    assign out[309] = in[594];
    assign out[540] = in[595];
    assign out[139] = in[596];
    assign out[3] = in[597];
    assign out[175] = in[598];
    assign out[471] = in[599];
    assign out[458] = in[600];
    assign out[617] = in[601];
    assign out[611] = in[602];
    assign out[430] = in[603];
    assign out[431] = in[604];
    assign out[274] = in[605];
    assign out[325] = in[606];
    assign out[200] = in[607];
    assign out[263] = in[608];
    assign out[186] = in[609];
    assign out[261] = in[610];
    assign out[326] = in[611];
    assign out[18] = in[612];
    assign out[76] = in[613];
    assign out[472] = in[614];
    assign out[330] = in[615];
    assign out[474] = in[616];
    assign out[193] = in[617];
    assign out[634] = in[618];
    assign out[13] = in[619];
    assign out[161] = in[620];
    assign out[521] = in[621];
    assign out[355] = in[622];
    assign out[639] = in[623];
    assign out[30] = in[624];
    assign out[22] = in[625];
    assign out[434] = in[626];
    assign out[591] = in[627];
    assign out[171] = in[628];
    assign out[362] = in[629];
    assign out[299] = in[630];
    assign out[575] = in[631];
    assign out[490] = in[632];
    assign out[176] = in[633];
    assign out[365] = in[634];
    assign out[515] = in[635];
    assign out[33] = in[636];
    assign out[415] = in[637];
    assign out[590] = in[638];
    assign out[497] = in[639];
endmodule

module odo_rotation_helper(in, out);
    input [63:0] in;
    output [63:0] out;
    assign out = {in[39:0], in[63:40]} ^ {in[58:0], in[63:59]} ^ {in[32:0], in[63:33]} ^ {in[30:0], in[63:31]} ^ {in[38:0], in[63:39]} ^ {in[46:0], in[63:47]};
endmodule

module odo_apply_rotations(in, out);
    input [639:0] in;
    output [639:0] out;
    wire [639:0] rot;
    odo_rotation_helper rot0inst(in[63:0], rot[63:0]);
    odo_rotation_helper rot1inst(in[127:64], rot[127:64]);
    odo_rotation_helper rot2inst(in[191:128], rot[191:128]);
    odo_rotation_helper rot3inst(in[255:192], rot[255:192]);
    odo_rotation_helper rot4inst(in[319:256], rot[319:256]);
    odo_rotation_helper rot5inst(in[383:320], rot[383:320]);
    odo_rotation_helper rot6inst(in[447:384], rot[447:384]);
    odo_rotation_helper rot7inst(in[511:448], rot[511:448]);
    odo_rotation_helper rot8inst(in[575:512], rot[575:512]);
    odo_rotation_helper rot9inst(in[639:576], rot[639:576]);
    assign out = rot ^ {in[63:0], in[639:64]};
endmodule

module odo_apply_round_key(key, in, out);
    input [9:0] key;
    input [639:0] in;
    output [639:0] out;
    assign out[0] = in[0] ^ key[0];
    assign out[63:1] = in[63:1];
    assign out[64] = in[64] ^ key[1];
    assign out[127:65] = in[127:65];
    assign out[128] = in[128] ^ key[2];
    assign out[191:129] = in[191:129];
    assign out[192] = in[192] ^ key[3];
    assign out[255:193] = in[255:193];
    assign out[256] = in[256] ^ key[4];
    assign out[319:257] = in[319:257];
    assign out[320] = in[320] ^ key[5];
    assign out[383:321] = in[383:321];
    assign out[384] = in[384] ^ key[6];
    assign out[447:385] = in[447:385];
    assign out[448] = in[448] ^ key[7];
    assign out[511:449] = in[511:449];
    assign out[512] = in[512] ^ key[8];
    assign out[575:513] = in[575:513];
    assign out[576] = in[576] ^ key[9];
    assign out[639:577] = in[639:577];
endmodule

module odo_full_round(clk, roundkey, in, out);
    input clk;
    input [9:0] roundkey;
    input [639:0] in;
    output [639:0] out;
    wire [639:0] mid[0:3];
    odo_apply_pbox0 pbox0inst(in, mid[0]);
    odo_apply_sboxes sboxes(clk, mid[0], mid[1]);
    odo_apply_pbox1 pbox1inst(mid[1], mid[2]);
    odo_apply_rotations rotations(mid[2], mid[3]);
    odo_apply_round_key keys(roundkey, mid[3], out);
endmodule

module odo_get_round_key0(clk, period, key);
    input clk;
    input [4:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        5'h00: key <= 10'h229;
        5'h01: key <= 10'h21d;
        5'h02: key <= 10'h006;
        5'h03: key <= 10'h07c;
        5'h04: key <= 10'h2f2;
        5'h05: key <= 10'h353;
        5'h06: key <= 10'h2f6;
        5'h07: key <= 10'h37f;
        5'h08: key <= 10'h029;
        5'h09: key <= 10'h153;
        5'h0a: key <= 10'h209;
        5'h0b: key <= 10'h3f3;
        5'h0c: key <= 10'h20e;
        5'h0d: key <= 10'h154;
        5'h0e: key <= 10'h1d6;
        5'h0f: key <= 10'h0f9;
        5'h10: key <= 10'h358;
        5'h11: key <= 10'h351;
        5'h12: key <= 10'h320;
        5'h13: key <= 10'h306;
        5'h14: key <= 10'h370;
    endcase
    end
endmodule

module odo_get_round_key1(clk, period, key);
    input clk;
    input [4:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        5'h00: key <= 10'h05a;
        5'h01: key <= 10'h3b6;
        5'h02: key <= 10'h3bb;
        5'h03: key <= 10'h0e8;
        5'h04: key <= 10'h35e;
        5'h05: key <= 10'h148;
        5'h06: key <= 10'h150;
        5'h07: key <= 10'h050;
        5'h08: key <= 10'h0e0;
        5'h09: key <= 10'h393;
        5'h0a: key <= 10'h1b0;
        5'h0b: key <= 10'h3c0;
        5'h0c: key <= 10'h158;
        5'h0d: key <= 10'h16e;
        5'h0e: key <= 10'h17c;
        5'h0f: key <= 10'h27e;
        5'h10: key <= 10'h17b;
        5'h11: key <= 10'h018;
        5'h12: key <= 10'h234;
        5'h13: key <= 10'h23d;
        5'h14: key <= 10'h0d2;
    endcase
    end
endmodule

module odo_get_round_key2(clk, period, key);
    input clk;
    input [4:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        5'h00: key <= 10'h3c9;
        5'h01: key <= 10'h2e0;
        5'h02: key <= 10'h26f;
        5'h03: key <= 10'h2b4;
        5'h04: key <= 10'h137;
        5'h05: key <= 10'h09b;
        5'h06: key <= 10'h17a;
        5'h07: key <= 10'h2fa;
        5'h08: key <= 10'h069;
        5'h09: key <= 10'h002;
        5'h0a: key <= 10'h1c4;
        5'h0b: key <= 10'h0fc;
        5'h0c: key <= 10'h089;
        5'h0d: key <= 10'h24e;
        5'h0e: key <= 10'h2be;
        5'h0f: key <= 10'h242;
        5'h10: key <= 10'h1cd;
        5'h11: key <= 10'h07e;
        5'h12: key <= 10'h1a0;
        5'h13: key <= 10'h09f;
        5'h14: key <= 10'h275;
    endcase
    end
endmodule

module odo_get_round_key3(clk, period, key);
    input clk;
    input [4:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        5'h00: key <= 10'h33f;
        5'h01: key <= 10'h3b8;
        5'h02: key <= 10'h0d3;
        5'h03: key <= 10'h078;
        5'h04: key <= 10'h3a0;
        5'h05: key <= 10'h07f;
        5'h06: key <= 10'h363;
        5'h07: key <= 10'h281;
        5'h08: key <= 10'h267;
        5'h09: key <= 10'h176;
        5'h0a: key <= 10'h0ec;
        5'h0b: key <= 10'h209;
        5'h0c: key <= 10'h1a4;
        5'h0d: key <= 10'h24e;
        5'h0e: key <= 10'h16d;
        5'h0f: key <= 10'h2df;
        5'h10: key <= 10'h169;
        5'h11: key <= 10'h0c2;
        5'h12: key <= 10'h125;
        5'h13: key <= 10'h061;
        5'h14: key <= 10'h227;
    endcase
    end
endmodule

module odo_encrypt_loop(clk, in, read, out, write);
    input clk;
    input [639:0] in;
    input read;
    output reg [639:0] out;
    output write;
    reg [639:0] state[3:0];
    wire [639:0] next[3:0];
    always @(posedge clk) state[1] <= next[0];
    always @(posedge clk) state[2] <= next[1];
    always @(posedge clk) state[3] <= next[2];
    wire [9:0] roundkey[3:0];
    reg [4:0] period[7:0];
    always @(posedge clk) period[1] <= period[0];
    always @(posedge clk) period[2] <= period[1];
    always @(posedge clk) period[3] <= period[2];
    always @(posedge clk) period[4] <= period[3];
    always @(posedge clk) period[5] <= period[4];
    always @(posedge clk) period[6] <= period[5];
    always @(posedge clk) period[7] <= period[6];
    odo_get_round_key0 get_key0(clk, period[0], roundkey[0]);
    odo_full_round round0(clk, roundkey[0], state[0], next[0]);
    odo_get_round_key1 get_key1(clk, period[2], roundkey[1]);
    odo_full_round round1(clk, roundkey[1], state[1], next[1]);
    odo_get_round_key2 get_key2(clk, period[4], roundkey[2]);
    odo_full_round round2(clk, roundkey[2], state[2], next[2]);
    odo_get_round_key3 get_key3(clk, period[6], roundkey[3]);
    odo_full_round round3(clk, roundkey[3], state[3], next[3]);
    always @(posedge clk) begin
        if (read)
        begin
            period[0] <= 0;
            state[0] <= in;
        end
        else
        begin
            period[0] <= period[7]+1;
            state[0] <= next[3];
        end
        out <= next[3];
    end
    reg [168:0] progress;
    initial progress = 169'h0;
    always @(posedge clk) progress[0] <= read;
    always @(posedge clk) progress[1] <= progress[0];
    always @(posedge clk) progress[2] <= progress[1];
    always @(posedge clk) progress[3] <= progress[2];
    always @(posedge clk) progress[4] <= progress[3];
    always @(posedge clk) progress[5] <= progress[4];
    always @(posedge clk) progress[6] <= progress[5];
    always @(posedge clk) progress[7] <= progress[6];
    always @(posedge clk) progress[8] <= progress[7];
    always @(posedge clk) progress[9] <= progress[8];
    always @(posedge clk) progress[10] <= progress[9];
    always @(posedge clk) progress[11] <= progress[10];
    always @(posedge clk) progress[12] <= progress[11];
    always @(posedge clk) progress[13] <= progress[12];
    always @(posedge clk) progress[14] <= progress[13];
    always @(posedge clk) progress[15] <= progress[14];
    always @(posedge clk) progress[16] <= progress[15];
    always @(posedge clk) progress[17] <= progress[16];
    always @(posedge clk) progress[18] <= progress[17];
    always @(posedge clk) progress[19] <= progress[18];
    always @(posedge clk) progress[20] <= progress[19];
    always @(posedge clk) progress[21] <= progress[20];
    always @(posedge clk) progress[22] <= progress[21];
    always @(posedge clk) progress[23] <= progress[22];
    always @(posedge clk) progress[24] <= progress[23];
    always @(posedge clk) progress[25] <= progress[24];
    always @(posedge clk) progress[26] <= progress[25];
    always @(posedge clk) progress[27] <= progress[26];
    always @(posedge clk) progress[28] <= progress[27];
    always @(posedge clk) progress[29] <= progress[28];
    always @(posedge clk) progress[30] <= progress[29];
    always @(posedge clk) progress[31] <= progress[30];
    always @(posedge clk) progress[32] <= progress[31];
    always @(posedge clk) progress[33] <= progress[32];
    always @(posedge clk) progress[34] <= progress[33];
    always @(posedge clk) progress[35] <= progress[34];
    always @(posedge clk) progress[36] <= progress[35];
    always @(posedge clk) progress[37] <= progress[36];
    always @(posedge clk) progress[38] <= progress[37];
    always @(posedge clk) progress[39] <= progress[38];
    always @(posedge clk) progress[40] <= progress[39];
    always @(posedge clk) progress[41] <= progress[40];
    always @(posedge clk) progress[42] <= progress[41];
    always @(posedge clk) progress[43] <= progress[42];
    always @(posedge clk) progress[44] <= progress[43];
    always @(posedge clk) progress[45] <= progress[44];
    always @(posedge clk) progress[46] <= progress[45];
    always @(posedge clk) progress[47] <= progress[46];
    always @(posedge clk) progress[48] <= progress[47];
    always @(posedge clk) progress[49] <= progress[48];
    always @(posedge clk) progress[50] <= progress[49];
    always @(posedge clk) progress[51] <= progress[50];
    always @(posedge clk) progress[52] <= progress[51];
    always @(posedge clk) progress[53] <= progress[52];
    always @(posedge clk) progress[54] <= progress[53];
    always @(posedge clk) progress[55] <= progress[54];
    always @(posedge clk) progress[56] <= progress[55];
    always @(posedge clk) progress[57] <= progress[56];
    always @(posedge clk) progress[58] <= progress[57];
    always @(posedge clk) progress[59] <= progress[58];
    always @(posedge clk) progress[60] <= progress[59];
    always @(posedge clk) progress[61] <= progress[60];
    always @(posedge clk) progress[62] <= progress[61];
    always @(posedge clk) progress[63] <= progress[62];
    always @(posedge clk) progress[64] <= progress[63];
    always @(posedge clk) progress[65] <= progress[64];
    always @(posedge clk) progress[66] <= progress[65];
    always @(posedge clk) progress[67] <= progress[66];
    always @(posedge clk) progress[68] <= progress[67];
    always @(posedge clk) progress[69] <= progress[68];
    always @(posedge clk) progress[70] <= progress[69];
    always @(posedge clk) progress[71] <= progress[70];
    always @(posedge clk) progress[72] <= progress[71];
    always @(posedge clk) progress[73] <= progress[72];
    always @(posedge clk) progress[74] <= progress[73];
    always @(posedge clk) progress[75] <= progress[74];
    always @(posedge clk) progress[76] <= progress[75];
    always @(posedge clk) progress[77] <= progress[76];
    always @(posedge clk) progress[78] <= progress[77];
    always @(posedge clk) progress[79] <= progress[78];
    always @(posedge clk) progress[80] <= progress[79];
    always @(posedge clk) progress[81] <= progress[80];
    always @(posedge clk) progress[82] <= progress[81];
    always @(posedge clk) progress[83] <= progress[82];
    always @(posedge clk) progress[84] <= progress[83];
    always @(posedge clk) progress[85] <= progress[84];
    always @(posedge clk) progress[86] <= progress[85];
    always @(posedge clk) progress[87] <= progress[86];
    always @(posedge clk) progress[88] <= progress[87];
    always @(posedge clk) progress[89] <= progress[88];
    always @(posedge clk) progress[90] <= progress[89];
    always @(posedge clk) progress[91] <= progress[90];
    always @(posedge clk) progress[92] <= progress[91];
    always @(posedge clk) progress[93] <= progress[92];
    always @(posedge clk) progress[94] <= progress[93];
    always @(posedge clk) progress[95] <= progress[94];
    always @(posedge clk) progress[96] <= progress[95];
    always @(posedge clk) progress[97] <= progress[96];
    always @(posedge clk) progress[98] <= progress[97];
    always @(posedge clk) progress[99] <= progress[98];
    always @(posedge clk) progress[100] <= progress[99];
    always @(posedge clk) progress[101] <= progress[100];
    always @(posedge clk) progress[102] <= progress[101];
    always @(posedge clk) progress[103] <= progress[102];
    always @(posedge clk) progress[104] <= progress[103];
    always @(posedge clk) progress[105] <= progress[104];
    always @(posedge clk) progress[106] <= progress[105];
    always @(posedge clk) progress[107] <= progress[106];
    always @(posedge clk) progress[108] <= progress[107];
    always @(posedge clk) progress[109] <= progress[108];
    always @(posedge clk) progress[110] <= progress[109];
    always @(posedge clk) progress[111] <= progress[110];
    always @(posedge clk) progress[112] <= progress[111];
    always @(posedge clk) progress[113] <= progress[112];
    always @(posedge clk) progress[114] <= progress[113];
    always @(posedge clk) progress[115] <= progress[114];
    always @(posedge clk) progress[116] <= progress[115];
    always @(posedge clk) progress[117] <= progress[116];
    always @(posedge clk) progress[118] <= progress[117];
    always @(posedge clk) progress[119] <= progress[118];
    always @(posedge clk) progress[120] <= progress[119];
    always @(posedge clk) progress[121] <= progress[120];
    always @(posedge clk) progress[122] <= progress[121];
    always @(posedge clk) progress[123] <= progress[122];
    always @(posedge clk) progress[124] <= progress[123];
    always @(posedge clk) progress[125] <= progress[124];
    always @(posedge clk) progress[126] <= progress[125];
    always @(posedge clk) progress[127] <= progress[126];
    always @(posedge clk) progress[128] <= progress[127];
    always @(posedge clk) progress[129] <= progress[128];
    always @(posedge clk) progress[130] <= progress[129];
    always @(posedge clk) progress[131] <= progress[130];
    always @(posedge clk) progress[132] <= progress[131];
    always @(posedge clk) progress[133] <= progress[132];
    always @(posedge clk) progress[134] <= progress[133];
    always @(posedge clk) progress[135] <= progress[134];
    always @(posedge clk) progress[136] <= progress[135];
    always @(posedge clk) progress[137] <= progress[136];
    always @(posedge clk) progress[138] <= progress[137];
    always @(posedge clk) progress[139] <= progress[138];
    always @(posedge clk) progress[140] <= progress[139];
    always @(posedge clk) progress[141] <= progress[140];
    always @(posedge clk) progress[142] <= progress[141];
    always @(posedge clk) progress[143] <= progress[142];
    always @(posedge clk) progress[144] <= progress[143];
    always @(posedge clk) progress[145] <= progress[144];
    always @(posedge clk) progress[146] <= progress[145];
    always @(posedge clk) progress[147] <= progress[146];
    always @(posedge clk) progress[148] <= progress[147];
    always @(posedge clk) progress[149] <= progress[148];
    always @(posedge clk) progress[150] <= progress[149];
    always @(posedge clk) progress[151] <= progress[150];
    always @(posedge clk) progress[152] <= progress[151];
    always @(posedge clk) progress[153] <= progress[152];
    always @(posedge clk) progress[154] <= progress[153];
    always @(posedge clk) progress[155] <= progress[154];
    always @(posedge clk) progress[156] <= progress[155];
    always @(posedge clk) progress[157] <= progress[156];
    always @(posedge clk) progress[158] <= progress[157];
    always @(posedge clk) progress[159] <= progress[158];
    always @(posedge clk) progress[160] <= progress[159];
    always @(posedge clk) progress[161] <= progress[160];
    always @(posedge clk) progress[162] <= progress[161];
    always @(posedge clk) progress[163] <= progress[162];
    always @(posedge clk) progress[164] <= progress[163];
    always @(posedge clk) progress[165] <= progress[164];
    always @(posedge clk) progress[166] <= progress[165];
    always @(posedge clk) progress[167] <= progress[166];
    always @(posedge clk) progress[168] <= progress[167];
    assign write = progress[168];
endmodule

module odo_encrypt(clk, in, read, out, write);
    localparam THROUGHPUT = 21;
    input clk;
    input [639:0] in;
    input read;
    output [639:0] out;
    output write;
    reg [1:0] progress;
    initial progress = 2'h0;
    reg [639:0] state[1:0];
    wire [639:0] next;
    odo_pre_mix premixer(state[0], next);
    odo_encrypt_loop crypter(clk, state[1], progress[1], out, write);
    always @(posedge clk) begin
        progress[0] <= read;
        progress[1] <= progress[0];
        state[0] <= in;
        state[1] <= next;
    end
endmodule